module c499_NOR_template (N1_PWL,N5_PWL,N9_PWL,N13_PWL,N17_PWL,N21_PWL,N25_PWL,N29_PWL,N33_PWL,N37_PWL,
            N41_PWL,N45_PWL,N49_PWL,N53_PWL,N57_PWL,N61_PWL,N65_PWL,N69_PWL,N73_PWL,N77_PWL,
            N81_PWL,N85_PWL,N89_PWL,N93_PWL,N97_PWL,N101_PWL,N105_PWL,N109_PWL,N113_PWL,N117_PWL,
            N121_PWL,N125_PWL,N129_PWL,N130_PWL,N131_PWL,N132_PWL,N133_PWL,N134_PWL,N135_PWL,N136_PWL,
            N137_PWL,N724_TERMINATION,N725_TERMINATION,N726_TERMINATION,N727_TERMINATION,N728_TERMINATION,
            N729_TERMINATION,N730_TERMINATION,N731_TERMINATION,N732_TERMINATION,N733_TERMINATION,
            N734_TERMINATION,N735_TERMINATION,N736_TERMINATION,N737_TERMINATION,N738_TERMINATION,
            N739_TERMINATION,N740_TERMINATION,N741_TERMINATION,N742_TERMINATION,N743_TERMINATION,
            N744_TERMINATION,N745_TERMINATION,N746_TERMINATION,N747_TERMINATION,N748_TERMINATION,
            N749_TERMINATION,N750_TERMINATION,N751_TERMINATION,N752_TERMINATION,N753_TERMINATION,
            N754_TERMINATION,N755_TERMINATION);

      input N1_PWL,N5_PWL,N9_PWL,N13_PWL,N17_PWL,N21_PWL,N25_PWL,N29_PWL,N33_PWL,N37_PWL,
            N41_PWL,N45_PWL,N49_PWL,N53_PWL,N57_PWL,N61_PWL,N65_PWL,N69_PWL,N73_PWL,N77_PWL,
            N81_PWL,N85_PWL,N89_PWL,N93_PWL,N97_PWL,N101_PWL,N105_PWL,N109_PWL,N113_PWL,N117_PWL,
            N121_PWL,N125_PWL,N129_PWL,N130_PWL,N131_PWL,N132_PWL,N133_PWL,N134_PWL,N135_PWL,N136_PWL,
            N137_PWL;

      output N724_TERMINATION,N725_TERMINATION,N726_TERMINATION,N727_TERMINATION,N728_TERMINATION,
            N729_TERMINATION,N730_TERMINATION,N731_TERMINATION,N732_TERMINATION,N733_TERMINATION,
            N734_TERMINATION,N735_TERMINATION,N736_TERMINATION,N737_TERMINATION,N738_TERMINATION,
            N739_TERMINATION,N740_TERMINATION,N741_TERMINATION,N742_TERMINATION,N743_TERMINATION,
            N744_TERMINATION,N745_TERMINATION,N746_TERMINATION,N747_TERMINATION,N748_TERMINATION,
            N749_TERMINATION,N750_TERMINATION,N751_TERMINATION,N752_TERMINATION,N753_TERMINATION,
            N754_TERMINATION,N755_TERMINATION;

      wire GND = 1'b0;
      wire XNOR_1_1_N1_PULSESHAPING_OUT, XNOR_1_2_N1_PULSESHAPING_OUT, XNOR_1_3_N1_PULSESHAPING_OUT, XNOR_1_4_N1_PULSESHAPING_OUT, XNOR_1_5_N1_PULSESHAPING_OUT, XNOR_1_6_N1_PULSESHAPING_OUT;
      NOR2_X1 XNOR_1_1_N1_PULSESHAPING (.ZN (XNOR_1_1_N1_PULSESHAPING_OUT), .A1 (N1_PWL), .A2 (GND));
      NOR2_X1 XNOR_1_2_N1_PULSESHAPING (.ZN (XNOR_1_2_N1_PULSESHAPING_OUT), .A1 (XNOR_1_1_N1_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_3_N1_PULSESHAPING (.ZN (XNOR_1_3_N1_PULSESHAPING_OUT), .A1 (XNOR_1_2_N1_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_4_N1_PULSESHAPING (.ZN (XNOR_1_4_N1_PULSESHAPING_OUT), .A1 (XNOR_1_3_N1_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_5_N1_PULSESHAPING (.ZN (XNOR_1_5_N1_PULSESHAPING_OUT), .A1 (XNOR_1_4_N1_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_6_N1_PULSESHAPING (.ZN (XNOR_1_6_N1_PULSESHAPING_OUT), .A1 (XNOR_1_5_N1_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_7_N1_PULSESHAPING (.ZN (N1), .A1 (XNOR_1_6_N1_PULSESHAPING_OUT), .A2 (GND));

      wire XNOR_1_1_N5_PULSESHAPING_OUT, XNOR_1_2_N5_PULSESHAPING_OUT, XNOR_1_3_N5_PULSESHAPING_OUT, XNOR_1_4_N5_PULSESHAPING_OUT, XNOR_1_5_N5_PULSESHAPING_OUT, XNOR_1_6_N5_PULSESHAPING_OUT;
      NOR2_X1 XNOR_1_1_N5_PULSESHAPING (.ZN (XNOR_1_1_N5_PULSESHAPING_OUT), .A1 (N5_PWL), .A2 (GND));
      NOR2_X1 XNOR_1_2_N5_PULSESHAPING (.ZN (XNOR_1_2_N5_PULSESHAPING_OUT), .A1 (XNOR_1_1_N5_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_3_N5_PULSESHAPING (.ZN (XNOR_1_3_N5_PULSESHAPING_OUT), .A1 (XNOR_1_2_N5_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_4_N5_PULSESHAPING (.ZN (XNOR_1_4_N5_PULSESHAPING_OUT), .A1 (XNOR_1_3_N5_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_5_N5_PULSESHAPING (.ZN (XNOR_1_5_N5_PULSESHAPING_OUT), .A1 (XNOR_1_4_N5_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_6_N5_PULSESHAPING (.ZN (XNOR_1_6_N5_PULSESHAPING_OUT), .A1 (XNOR_1_5_N5_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_7_N5_PULSESHAPING (.ZN (N5), .A1 (XNOR_1_6_N5_PULSESHAPING_OUT), .A2 (GND));

      wire XNOR_1_1_N9_PULSESHAPING_OUT, XNOR_1_2_N9_PULSESHAPING_OUT, XNOR_1_3_N9_PULSESHAPING_OUT, XNOR_1_4_N9_PULSESHAPING_OUT, XNOR_1_5_N9_PULSESHAPING_OUT, XNOR_1_6_N9_PULSESHAPING_OUT;
      NOR2_X1 XNOR_1_1_N9_PULSESHAPING (.ZN (XNOR_1_1_N9_PULSESHAPING_OUT), .A1 (N9_PWL), .A2 (GND));
      NOR2_X1 XNOR_1_2_N9_PULSESHAPING (.ZN (XNOR_1_2_N9_PULSESHAPING_OUT), .A1 (XNOR_1_1_N9_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_3_N9_PULSESHAPING (.ZN (XNOR_1_3_N9_PULSESHAPING_OUT), .A1 (XNOR_1_2_N9_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_4_N9_PULSESHAPING (.ZN (XNOR_1_4_N9_PULSESHAPING_OUT), .A1 (XNOR_1_3_N9_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_5_N9_PULSESHAPING (.ZN (XNOR_1_5_N9_PULSESHAPING_OUT), .A1 (XNOR_1_4_N9_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_6_N9_PULSESHAPING (.ZN (XNOR_1_6_N9_PULSESHAPING_OUT), .A1 (XNOR_1_5_N9_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_7_N9_PULSESHAPING (.ZN (N9), .A1 (XNOR_1_6_N9_PULSESHAPING_OUT), .A2 (GND));

      wire XNOR_1_1_N13_PULSESHAPING_OUT, XNOR_1_2_N13_PULSESHAPING_OUT, XNOR_1_3_N13_PULSESHAPING_OUT, XNOR_1_4_N13_PULSESHAPING_OUT, XNOR_1_5_N13_PULSESHAPING_OUT, XNOR_1_6_N13_PULSESHAPING_OUT;
      NOR2_X1 XNOR_1_1_N13_PULSESHAPING (.ZN (XNOR_1_1_N13_PULSESHAPING_OUT), .A1 (N13_PWL), .A2 (GND));
      NOR2_X1 XNOR_1_2_N13_PULSESHAPING (.ZN (XNOR_1_2_N13_PULSESHAPING_OUT), .A1 (XNOR_1_1_N13_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_3_N13_PULSESHAPING (.ZN (XNOR_1_3_N13_PULSESHAPING_OUT), .A1 (XNOR_1_2_N13_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_4_N13_PULSESHAPING (.ZN (XNOR_1_4_N13_PULSESHAPING_OUT), .A1 (XNOR_1_3_N13_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_5_N13_PULSESHAPING (.ZN (XNOR_1_5_N13_PULSESHAPING_OUT), .A1 (XNOR_1_4_N13_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_6_N13_PULSESHAPING (.ZN (XNOR_1_6_N13_PULSESHAPING_OUT), .A1 (XNOR_1_5_N13_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_7_N13_PULSESHAPING (.ZN (N13), .A1 (XNOR_1_6_N13_PULSESHAPING_OUT), .A2 (GND));

      wire XNOR_1_1_N17_PULSESHAPING_OUT, XNOR_1_2_N17_PULSESHAPING_OUT, XNOR_1_3_N17_PULSESHAPING_OUT, XNOR_1_4_N17_PULSESHAPING_OUT, XNOR_1_5_N17_PULSESHAPING_OUT, XNOR_1_6_N17_PULSESHAPING_OUT;
      NOR2_X1 XNOR_1_1_N17_PULSESHAPING (.ZN (XNOR_1_1_N17_PULSESHAPING_OUT), .A1 (N17_PWL), .A2 (GND));
      NOR2_X1 XNOR_1_2_N17_PULSESHAPING (.ZN (XNOR_1_2_N17_PULSESHAPING_OUT), .A1 (XNOR_1_1_N17_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_3_N17_PULSESHAPING (.ZN (XNOR_1_3_N17_PULSESHAPING_OUT), .A1 (XNOR_1_2_N17_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_4_N17_PULSESHAPING (.ZN (XNOR_1_4_N17_PULSESHAPING_OUT), .A1 (XNOR_1_3_N17_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_5_N17_PULSESHAPING (.ZN (XNOR_1_5_N17_PULSESHAPING_OUT), .A1 (XNOR_1_4_N17_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_6_N17_PULSESHAPING (.ZN (XNOR_1_6_N17_PULSESHAPING_OUT), .A1 (XNOR_1_5_N17_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_7_N17_PULSESHAPING (.ZN (N17), .A1 (XNOR_1_6_N17_PULSESHAPING_OUT), .A2 (GND));

      wire XNOR_1_1_N21_PULSESHAPING_OUT, XNOR_1_2_N21_PULSESHAPING_OUT, XNOR_1_3_N21_PULSESHAPING_OUT, XNOR_1_4_N21_PULSESHAPING_OUT, XNOR_1_5_N21_PULSESHAPING_OUT, XNOR_1_6_N21_PULSESHAPING_OUT;
      NOR2_X1 XNOR_1_1_N21_PULSESHAPING (.ZN (XNOR_1_1_N21_PULSESHAPING_OUT), .A1 (N21_PWL), .A2 (GND));
      NOR2_X1 XNOR_1_2_N21_PULSESHAPING (.ZN (XNOR_1_2_N21_PULSESHAPING_OUT), .A1 (XNOR_1_1_N21_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_3_N21_PULSESHAPING (.ZN (XNOR_1_3_N21_PULSESHAPING_OUT), .A1 (XNOR_1_2_N21_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_4_N21_PULSESHAPING (.ZN (XNOR_1_4_N21_PULSESHAPING_OUT), .A1 (XNOR_1_3_N21_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_5_N21_PULSESHAPING (.ZN (XNOR_1_5_N21_PULSESHAPING_OUT), .A1 (XNOR_1_4_N21_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_6_N21_PULSESHAPING (.ZN (XNOR_1_6_N21_PULSESHAPING_OUT), .A1 (XNOR_1_5_N21_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_7_N21_PULSESHAPING (.ZN (N21), .A1 (XNOR_1_6_N21_PULSESHAPING_OUT), .A2 (GND));

      wire XNOR_1_1_N25_PULSESHAPING_OUT, XNOR_1_2_N25_PULSESHAPING_OUT, XNOR_1_3_N25_PULSESHAPING_OUT, XNOR_1_4_N25_PULSESHAPING_OUT, XNOR_1_5_N25_PULSESHAPING_OUT, XNOR_1_6_N25_PULSESHAPING_OUT;
      NOR2_X1 XNOR_1_1_N25_PULSESHAPING (.ZN (XNOR_1_1_N25_PULSESHAPING_OUT), .A1 (N25_PWL), .A2 (GND));
      NOR2_X1 XNOR_1_2_N25_PULSESHAPING (.ZN (XNOR_1_2_N25_PULSESHAPING_OUT), .A1 (XNOR_1_1_N25_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_3_N25_PULSESHAPING (.ZN (XNOR_1_3_N25_PULSESHAPING_OUT), .A1 (XNOR_1_2_N25_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_4_N25_PULSESHAPING (.ZN (XNOR_1_4_N25_PULSESHAPING_OUT), .A1 (XNOR_1_3_N25_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_5_N25_PULSESHAPING (.ZN (XNOR_1_5_N25_PULSESHAPING_OUT), .A1 (XNOR_1_4_N25_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_6_N25_PULSESHAPING (.ZN (XNOR_1_6_N25_PULSESHAPING_OUT), .A1 (XNOR_1_5_N25_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_7_N25_PULSESHAPING (.ZN (N25), .A1 (XNOR_1_6_N25_PULSESHAPING_OUT), .A2 (GND));

      wire XNOR_1_1_N29_PULSESHAPING_OUT, XNOR_1_2_N29_PULSESHAPING_OUT, XNOR_1_3_N29_PULSESHAPING_OUT, XNOR_1_4_N29_PULSESHAPING_OUT, XNOR_1_5_N29_PULSESHAPING_OUT, XNOR_1_6_N29_PULSESHAPING_OUT;
      NOR2_X1 XNOR_1_1_N29_PULSESHAPING (.ZN (XNOR_1_1_N29_PULSESHAPING_OUT), .A1 (N29_PWL), .A2 (GND));
      NOR2_X1 XNOR_1_2_N29_PULSESHAPING (.ZN (XNOR_1_2_N29_PULSESHAPING_OUT), .A1 (XNOR_1_1_N29_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_3_N29_PULSESHAPING (.ZN (XNOR_1_3_N29_PULSESHAPING_OUT), .A1 (XNOR_1_2_N29_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_4_N29_PULSESHAPING (.ZN (XNOR_1_4_N29_PULSESHAPING_OUT), .A1 (XNOR_1_3_N29_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_5_N29_PULSESHAPING (.ZN (XNOR_1_5_N29_PULSESHAPING_OUT), .A1 (XNOR_1_4_N29_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_6_N29_PULSESHAPING (.ZN (XNOR_1_6_N29_PULSESHAPING_OUT), .A1 (XNOR_1_5_N29_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_7_N29_PULSESHAPING (.ZN (N29), .A1 (XNOR_1_6_N29_PULSESHAPING_OUT), .A2 (GND));

      wire XNOR_1_1_N33_PULSESHAPING_OUT, XNOR_1_2_N33_PULSESHAPING_OUT, XNOR_1_3_N33_PULSESHAPING_OUT, XNOR_1_4_N33_PULSESHAPING_OUT, XNOR_1_5_N33_PULSESHAPING_OUT, XNOR_1_6_N33_PULSESHAPING_OUT;
      NOR2_X1 XNOR_1_1_N33_PULSESHAPING (.ZN (XNOR_1_1_N33_PULSESHAPING_OUT), .A1 (N33_PWL), .A2 (GND));
      NOR2_X1 XNOR_1_2_N33_PULSESHAPING (.ZN (XNOR_1_2_N33_PULSESHAPING_OUT), .A1 (XNOR_1_1_N33_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_3_N33_PULSESHAPING (.ZN (XNOR_1_3_N33_PULSESHAPING_OUT), .A1 (XNOR_1_2_N33_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_4_N33_PULSESHAPING (.ZN (XNOR_1_4_N33_PULSESHAPING_OUT), .A1 (XNOR_1_3_N33_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_5_N33_PULSESHAPING (.ZN (XNOR_1_5_N33_PULSESHAPING_OUT), .A1 (XNOR_1_4_N33_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_6_N33_PULSESHAPING (.ZN (XNOR_1_6_N33_PULSESHAPING_OUT), .A1 (XNOR_1_5_N33_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_7_N33_PULSESHAPING (.ZN (N33), .A1 (XNOR_1_6_N33_PULSESHAPING_OUT), .A2 (GND));

      wire XNOR_1_1_N37_PULSESHAPING_OUT, XNOR_1_2_N37_PULSESHAPING_OUT, XNOR_1_3_N37_PULSESHAPING_OUT, XNOR_1_4_N37_PULSESHAPING_OUT, XNOR_1_5_N37_PULSESHAPING_OUT, XNOR_1_6_N37_PULSESHAPING_OUT;
      NOR2_X1 XNOR_1_1_N37_PULSESHAPING (.ZN (XNOR_1_1_N37_PULSESHAPING_OUT), .A1 (N37_PWL), .A2 (GND));
      NOR2_X1 XNOR_1_2_N37_PULSESHAPING (.ZN (XNOR_1_2_N37_PULSESHAPING_OUT), .A1 (XNOR_1_1_N37_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_3_N37_PULSESHAPING (.ZN (XNOR_1_3_N37_PULSESHAPING_OUT), .A1 (XNOR_1_2_N37_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_4_N37_PULSESHAPING (.ZN (XNOR_1_4_N37_PULSESHAPING_OUT), .A1 (XNOR_1_3_N37_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_5_N37_PULSESHAPING (.ZN (XNOR_1_5_N37_PULSESHAPING_OUT), .A1 (XNOR_1_4_N37_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_6_N37_PULSESHAPING (.ZN (XNOR_1_6_N37_PULSESHAPING_OUT), .A1 (XNOR_1_5_N37_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_7_N37_PULSESHAPING (.ZN (N37), .A1 (XNOR_1_6_N37_PULSESHAPING_OUT), .A2 (GND));

      wire XNOR_1_1_N41_PULSESHAPING_OUT, XNOR_1_2_N41_PULSESHAPING_OUT, XNOR_1_3_N41_PULSESHAPING_OUT, XNOR_1_4_N41_PULSESHAPING_OUT, XNOR_1_5_N41_PULSESHAPING_OUT, XNOR_1_6_N41_PULSESHAPING_OUT;
      NOR2_X1 XNOR_1_1_N41_PULSESHAPING (.ZN (XNOR_1_1_N41_PULSESHAPING_OUT), .A1 (N41_PWL), .A2 (GND));
      NOR2_X1 XNOR_1_2_N41_PULSESHAPING (.ZN (XNOR_1_2_N41_PULSESHAPING_OUT), .A1 (XNOR_1_1_N41_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_3_N41_PULSESHAPING (.ZN (XNOR_1_3_N41_PULSESHAPING_OUT), .A1 (XNOR_1_2_N41_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_4_N41_PULSESHAPING (.ZN (XNOR_1_4_N41_PULSESHAPING_OUT), .A1 (XNOR_1_3_N41_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_5_N41_PULSESHAPING (.ZN (XNOR_1_5_N41_PULSESHAPING_OUT), .A1 (XNOR_1_4_N41_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_6_N41_PULSESHAPING (.ZN (XNOR_1_6_N41_PULSESHAPING_OUT), .A1 (XNOR_1_5_N41_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_7_N41_PULSESHAPING (.ZN (N41), .A1 (XNOR_1_6_N41_PULSESHAPING_OUT), .A2 (GND));

      wire XNOR_1_1_N45_PULSESHAPING_OUT, XNOR_1_2_N45_PULSESHAPING_OUT, XNOR_1_3_N45_PULSESHAPING_OUT, XNOR_1_4_N45_PULSESHAPING_OUT, XNOR_1_5_N45_PULSESHAPING_OUT, XNOR_1_6_N45_PULSESHAPING_OUT;
      NOR2_X1 XNOR_1_1_N45_PULSESHAPING (.ZN (XNOR_1_1_N45_PULSESHAPING_OUT), .A1 (N45_PWL), .A2 (GND));
      NOR2_X1 XNOR_1_2_N45_PULSESHAPING (.ZN (XNOR_1_2_N45_PULSESHAPING_OUT), .A1 (XNOR_1_1_N45_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_3_N45_PULSESHAPING (.ZN (XNOR_1_3_N45_PULSESHAPING_OUT), .A1 (XNOR_1_2_N45_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_4_N45_PULSESHAPING (.ZN (XNOR_1_4_N45_PULSESHAPING_OUT), .A1 (XNOR_1_3_N45_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_5_N45_PULSESHAPING (.ZN (XNOR_1_5_N45_PULSESHAPING_OUT), .A1 (XNOR_1_4_N45_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_6_N45_PULSESHAPING (.ZN (XNOR_1_6_N45_PULSESHAPING_OUT), .A1 (XNOR_1_5_N45_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_7_N45_PULSESHAPING (.ZN (N45), .A1 (XNOR_1_6_N45_PULSESHAPING_OUT), .A2 (GND));

      wire XNOR_1_1_N49_PULSESHAPING_OUT, XNOR_1_2_N49_PULSESHAPING_OUT, XNOR_1_3_N49_PULSESHAPING_OUT, XNOR_1_4_N49_PULSESHAPING_OUT, XNOR_1_5_N49_PULSESHAPING_OUT, XNOR_1_6_N49_PULSESHAPING_OUT;
      NOR2_X1 XNOR_1_1_N49_PULSESHAPING (.ZN (XNOR_1_1_N49_PULSESHAPING_OUT), .A1 (N49_PWL), .A2 (GND));
      NOR2_X1 XNOR_1_2_N49_PULSESHAPING (.ZN (XNOR_1_2_N49_PULSESHAPING_OUT), .A1 (XNOR_1_1_N49_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_3_N49_PULSESHAPING (.ZN (XNOR_1_3_N49_PULSESHAPING_OUT), .A1 (XNOR_1_2_N49_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_4_N49_PULSESHAPING (.ZN (XNOR_1_4_N49_PULSESHAPING_OUT), .A1 (XNOR_1_3_N49_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_5_N49_PULSESHAPING (.ZN (XNOR_1_5_N49_PULSESHAPING_OUT), .A1 (XNOR_1_4_N49_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_6_N49_PULSESHAPING (.ZN (XNOR_1_6_N49_PULSESHAPING_OUT), .A1 (XNOR_1_5_N49_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_7_N49_PULSESHAPING (.ZN (N49), .A1 (XNOR_1_6_N49_PULSESHAPING_OUT), .A2 (GND));

      wire XNOR_1_1_N53_PULSESHAPING_OUT, XNOR_1_2_N53_PULSESHAPING_OUT, XNOR_1_3_N53_PULSESHAPING_OUT, XNOR_1_4_N53_PULSESHAPING_OUT, XNOR_1_5_N53_PULSESHAPING_OUT, XNOR_1_6_N53_PULSESHAPING_OUT;
      NOR2_X1 XNOR_1_1_N53_PULSESHAPING (.ZN (XNOR_1_1_N53_PULSESHAPING_OUT), .A1 (N53_PWL), .A2 (GND));
      NOR2_X1 XNOR_1_2_N53_PULSESHAPING (.ZN (XNOR_1_2_N53_PULSESHAPING_OUT), .A1 (XNOR_1_1_N53_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_3_N53_PULSESHAPING (.ZN (XNOR_1_3_N53_PULSESHAPING_OUT), .A1 (XNOR_1_2_N53_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_4_N53_PULSESHAPING (.ZN (XNOR_1_4_N53_PULSESHAPING_OUT), .A1 (XNOR_1_3_N53_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_5_N53_PULSESHAPING (.ZN (XNOR_1_5_N53_PULSESHAPING_OUT), .A1 (XNOR_1_4_N53_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_6_N53_PULSESHAPING (.ZN (XNOR_1_6_N53_PULSESHAPING_OUT), .A1 (XNOR_1_5_N53_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_7_N53_PULSESHAPING (.ZN (N53), .A1 (XNOR_1_6_N53_PULSESHAPING_OUT), .A2 (GND));

      wire XNOR_1_1_N57_PULSESHAPING_OUT, XNOR_1_2_N57_PULSESHAPING_OUT, XNOR_1_3_N57_PULSESHAPING_OUT, XNOR_1_4_N57_PULSESHAPING_OUT, XNOR_1_5_N57_PULSESHAPING_OUT, XNOR_1_6_N57_PULSESHAPING_OUT;
      NOR2_X1 XNOR_1_1_N57_PULSESHAPING (.ZN (XNOR_1_1_N57_PULSESHAPING_OUT), .A1 (N57_PWL), .A2 (GND));
      NOR2_X1 XNOR_1_2_N57_PULSESHAPING (.ZN (XNOR_1_2_N57_PULSESHAPING_OUT), .A1 (XNOR_1_1_N57_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_3_N57_PULSESHAPING (.ZN (XNOR_1_3_N57_PULSESHAPING_OUT), .A1 (XNOR_1_2_N57_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_4_N57_PULSESHAPING (.ZN (XNOR_1_4_N57_PULSESHAPING_OUT), .A1 (XNOR_1_3_N57_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_5_N57_PULSESHAPING (.ZN (XNOR_1_5_N57_PULSESHAPING_OUT), .A1 (XNOR_1_4_N57_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_6_N57_PULSESHAPING (.ZN (XNOR_1_6_N57_PULSESHAPING_OUT), .A1 (XNOR_1_5_N57_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_7_N57_PULSESHAPING (.ZN (N57), .A1 (XNOR_1_6_N57_PULSESHAPING_OUT), .A2 (GND));

      wire XNOR_1_1_N61_PULSESHAPING_OUT, XNOR_1_2_N61_PULSESHAPING_OUT, XNOR_1_3_N61_PULSESHAPING_OUT, XNOR_1_4_N61_PULSESHAPING_OUT, XNOR_1_5_N61_PULSESHAPING_OUT, XNOR_1_6_N61_PULSESHAPING_OUT;
      NOR2_X1 XNOR_1_1_N61_PULSESHAPING (.ZN (XNOR_1_1_N61_PULSESHAPING_OUT), .A1 (N61_PWL), .A2 (GND));
      NOR2_X1 XNOR_1_2_N61_PULSESHAPING (.ZN (XNOR_1_2_N61_PULSESHAPING_OUT), .A1 (XNOR_1_1_N61_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_3_N61_PULSESHAPING (.ZN (XNOR_1_3_N61_PULSESHAPING_OUT), .A1 (XNOR_1_2_N61_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_4_N61_PULSESHAPING (.ZN (XNOR_1_4_N61_PULSESHAPING_OUT), .A1 (XNOR_1_3_N61_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_5_N61_PULSESHAPING (.ZN (XNOR_1_5_N61_PULSESHAPING_OUT), .A1 (XNOR_1_4_N61_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_6_N61_PULSESHAPING (.ZN (XNOR_1_6_N61_PULSESHAPING_OUT), .A1 (XNOR_1_5_N61_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_7_N61_PULSESHAPING (.ZN (N61), .A1 (XNOR_1_6_N61_PULSESHAPING_OUT), .A2 (GND));

      wire XNOR_1_1_N65_PULSESHAPING_OUT, XNOR_1_2_N65_PULSESHAPING_OUT, XNOR_1_3_N65_PULSESHAPING_OUT, XNOR_1_4_N65_PULSESHAPING_OUT, XNOR_1_5_N65_PULSESHAPING_OUT, XNOR_1_6_N65_PULSESHAPING_OUT;
      NOR2_X1 XNOR_1_1_N65_PULSESHAPING (.ZN (XNOR_1_1_N65_PULSESHAPING_OUT), .A1 (N65_PWL), .A2 (GND));
      NOR2_X1 XNOR_1_2_N65_PULSESHAPING (.ZN (XNOR_1_2_N65_PULSESHAPING_OUT), .A1 (XNOR_1_1_N65_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_3_N65_PULSESHAPING (.ZN (XNOR_1_3_N65_PULSESHAPING_OUT), .A1 (XNOR_1_2_N65_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_4_N65_PULSESHAPING (.ZN (XNOR_1_4_N65_PULSESHAPING_OUT), .A1 (XNOR_1_3_N65_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_5_N65_PULSESHAPING (.ZN (XNOR_1_5_N65_PULSESHAPING_OUT), .A1 (XNOR_1_4_N65_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_6_N65_PULSESHAPING (.ZN (XNOR_1_6_N65_PULSESHAPING_OUT), .A1 (XNOR_1_5_N65_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_7_N65_PULSESHAPING (.ZN (N65), .A1 (XNOR_1_6_N65_PULSESHAPING_OUT), .A2 (GND));

      wire XNOR_1_1_N69_PULSESHAPING_OUT, XNOR_1_2_N69_PULSESHAPING_OUT, XNOR_1_3_N69_PULSESHAPING_OUT, XNOR_1_4_N69_PULSESHAPING_OUT, XNOR_1_5_N69_PULSESHAPING_OUT, XNOR_1_6_N69_PULSESHAPING_OUT;
      NOR2_X1 XNOR_1_1_N69_PULSESHAPING (.ZN (XNOR_1_1_N69_PULSESHAPING_OUT), .A1 (N69_PWL), .A2 (GND));
      NOR2_X1 XNOR_1_2_N69_PULSESHAPING (.ZN (XNOR_1_2_N69_PULSESHAPING_OUT), .A1 (XNOR_1_1_N69_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_3_N69_PULSESHAPING (.ZN (XNOR_1_3_N69_PULSESHAPING_OUT), .A1 (XNOR_1_2_N69_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_4_N69_PULSESHAPING (.ZN (XNOR_1_4_N69_PULSESHAPING_OUT), .A1 (XNOR_1_3_N69_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_5_N69_PULSESHAPING (.ZN (XNOR_1_5_N69_PULSESHAPING_OUT), .A1 (XNOR_1_4_N69_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_6_N69_PULSESHAPING (.ZN (XNOR_1_6_N69_PULSESHAPING_OUT), .A1 (XNOR_1_5_N69_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_7_N69_PULSESHAPING (.ZN (N69), .A1 (XNOR_1_6_N69_PULSESHAPING_OUT), .A2 (GND));

      wire XNOR_1_1_N73_PULSESHAPING_OUT, XNOR_1_2_N73_PULSESHAPING_OUT, XNOR_1_3_N73_PULSESHAPING_OUT, XNOR_1_4_N73_PULSESHAPING_OUT, XNOR_1_5_N73_PULSESHAPING_OUT, XNOR_1_6_N73_PULSESHAPING_OUT;
      NOR2_X1 XNOR_1_1_N73_PULSESHAPING (.ZN (XNOR_1_1_N73_PULSESHAPING_OUT), .A1 (N73_PWL), .A2 (GND));
      NOR2_X1 XNOR_1_2_N73_PULSESHAPING (.ZN (XNOR_1_2_N73_PULSESHAPING_OUT), .A1 (XNOR_1_1_N73_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_3_N73_PULSESHAPING (.ZN (XNOR_1_3_N73_PULSESHAPING_OUT), .A1 (XNOR_1_2_N73_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_4_N73_PULSESHAPING (.ZN (XNOR_1_4_N73_PULSESHAPING_OUT), .A1 (XNOR_1_3_N73_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_5_N73_PULSESHAPING (.ZN (XNOR_1_5_N73_PULSESHAPING_OUT), .A1 (XNOR_1_4_N73_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_6_N73_PULSESHAPING (.ZN (XNOR_1_6_N73_PULSESHAPING_OUT), .A1 (XNOR_1_5_N73_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_7_N73_PULSESHAPING (.ZN (N73), .A1 (XNOR_1_6_N73_PULSESHAPING_OUT), .A2 (GND));

      wire XNOR_1_1_N77_PULSESHAPING_OUT, XNOR_1_2_N77_PULSESHAPING_OUT, XNOR_1_3_N77_PULSESHAPING_OUT, XNOR_1_4_N77_PULSESHAPING_OUT, XNOR_1_5_N77_PULSESHAPING_OUT, XNOR_1_6_N77_PULSESHAPING_OUT;
      NOR2_X1 XNOR_1_1_N77_PULSESHAPING (.ZN (XNOR_1_1_N77_PULSESHAPING_OUT), .A1 (N77_PWL), .A2 (GND));
      NOR2_X1 XNOR_1_2_N77_PULSESHAPING (.ZN (XNOR_1_2_N77_PULSESHAPING_OUT), .A1 (XNOR_1_1_N77_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_3_N77_PULSESHAPING (.ZN (XNOR_1_3_N77_PULSESHAPING_OUT), .A1 (XNOR_1_2_N77_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_4_N77_PULSESHAPING (.ZN (XNOR_1_4_N77_PULSESHAPING_OUT), .A1 (XNOR_1_3_N77_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_5_N77_PULSESHAPING (.ZN (XNOR_1_5_N77_PULSESHAPING_OUT), .A1 (XNOR_1_4_N77_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_6_N77_PULSESHAPING (.ZN (XNOR_1_6_N77_PULSESHAPING_OUT), .A1 (XNOR_1_5_N77_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_7_N77_PULSESHAPING (.ZN (N77), .A1 (XNOR_1_6_N77_PULSESHAPING_OUT), .A2 (GND));

      wire XNOR_1_1_N81_PULSESHAPING_OUT, XNOR_1_2_N81_PULSESHAPING_OUT, XNOR_1_3_N81_PULSESHAPING_OUT, XNOR_1_4_N81_PULSESHAPING_OUT, XNOR_1_5_N81_PULSESHAPING_OUT, XNOR_1_6_N81_PULSESHAPING_OUT;
      NOR2_X1 XNOR_1_1_N81_PULSESHAPING (.ZN (XNOR_1_1_N81_PULSESHAPING_OUT), .A1 (N81_PWL), .A2 (GND));
      NOR2_X1 XNOR_1_2_N81_PULSESHAPING (.ZN (XNOR_1_2_N81_PULSESHAPING_OUT), .A1 (XNOR_1_1_N81_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_3_N81_PULSESHAPING (.ZN (XNOR_1_3_N81_PULSESHAPING_OUT), .A1 (XNOR_1_2_N81_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_4_N81_PULSESHAPING (.ZN (XNOR_1_4_N81_PULSESHAPING_OUT), .A1 (XNOR_1_3_N81_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_5_N81_PULSESHAPING (.ZN (XNOR_1_5_N81_PULSESHAPING_OUT), .A1 (XNOR_1_4_N81_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_6_N81_PULSESHAPING (.ZN (XNOR_1_6_N81_PULSESHAPING_OUT), .A1 (XNOR_1_5_N81_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_7_N81_PULSESHAPING (.ZN (N81), .A1 (XNOR_1_6_N81_PULSESHAPING_OUT), .A2 (GND));

      wire XNOR_1_1_N85_PULSESHAPING_OUT, XNOR_1_2_N85_PULSESHAPING_OUT, XNOR_1_3_N85_PULSESHAPING_OUT, XNOR_1_4_N85_PULSESHAPING_OUT, XNOR_1_5_N85_PULSESHAPING_OUT, XNOR_1_6_N85_PULSESHAPING_OUT;
      NOR2_X1 XNOR_1_1_N85_PULSESHAPING (.ZN (XNOR_1_1_N85_PULSESHAPING_OUT), .A1 (N85_PWL), .A2 (GND));
      NOR2_X1 XNOR_1_2_N85_PULSESHAPING (.ZN (XNOR_1_2_N85_PULSESHAPING_OUT), .A1 (XNOR_1_1_N85_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_3_N85_PULSESHAPING (.ZN (XNOR_1_3_N85_PULSESHAPING_OUT), .A1 (XNOR_1_2_N85_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_4_N85_PULSESHAPING (.ZN (XNOR_1_4_N85_PULSESHAPING_OUT), .A1 (XNOR_1_3_N85_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_5_N85_PULSESHAPING (.ZN (XNOR_1_5_N85_PULSESHAPING_OUT), .A1 (XNOR_1_4_N85_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_6_N85_PULSESHAPING (.ZN (XNOR_1_6_N85_PULSESHAPING_OUT), .A1 (XNOR_1_5_N85_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_7_N85_PULSESHAPING (.ZN (N85), .A1 (XNOR_1_6_N85_PULSESHAPING_OUT), .A2 (GND));

      wire XNOR_1_1_N89_PULSESHAPING_OUT, XNOR_1_2_N89_PULSESHAPING_OUT, XNOR_1_3_N89_PULSESHAPING_OUT, XNOR_1_4_N89_PULSESHAPING_OUT, XNOR_1_5_N89_PULSESHAPING_OUT, XNOR_1_6_N89_PULSESHAPING_OUT;
      NOR2_X1 XNOR_1_1_N89_PULSESHAPING (.ZN (XNOR_1_1_N89_PULSESHAPING_OUT), .A1 (N89_PWL), .A2 (GND));
      NOR2_X1 XNOR_1_2_N89_PULSESHAPING (.ZN (XNOR_1_2_N89_PULSESHAPING_OUT), .A1 (XNOR_1_1_N89_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_3_N89_PULSESHAPING (.ZN (XNOR_1_3_N89_PULSESHAPING_OUT), .A1 (XNOR_1_2_N89_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_4_N89_PULSESHAPING (.ZN (XNOR_1_4_N89_PULSESHAPING_OUT), .A1 (XNOR_1_3_N89_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_5_N89_PULSESHAPING (.ZN (XNOR_1_5_N89_PULSESHAPING_OUT), .A1 (XNOR_1_4_N89_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_6_N89_PULSESHAPING (.ZN (XNOR_1_6_N89_PULSESHAPING_OUT), .A1 (XNOR_1_5_N89_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_7_N89_PULSESHAPING (.ZN (N89), .A1 (XNOR_1_6_N89_PULSESHAPING_OUT), .A2 (GND));

      wire XNOR_1_1_N93_PULSESHAPING_OUT, XNOR_1_2_N93_PULSESHAPING_OUT, XNOR_1_3_N93_PULSESHAPING_OUT, XNOR_1_4_N93_PULSESHAPING_OUT, XNOR_1_5_N93_PULSESHAPING_OUT, XNOR_1_6_N93_PULSESHAPING_OUT;
      NOR2_X1 XNOR_1_1_N93_PULSESHAPING (.ZN (XNOR_1_1_N93_PULSESHAPING_OUT), .A1 (N93_PWL), .A2 (GND));
      NOR2_X1 XNOR_1_2_N93_PULSESHAPING (.ZN (XNOR_1_2_N93_PULSESHAPING_OUT), .A1 (XNOR_1_1_N93_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_3_N93_PULSESHAPING (.ZN (XNOR_1_3_N93_PULSESHAPING_OUT), .A1 (XNOR_1_2_N93_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_4_N93_PULSESHAPING (.ZN (XNOR_1_4_N93_PULSESHAPING_OUT), .A1 (XNOR_1_3_N93_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_5_N93_PULSESHAPING (.ZN (XNOR_1_5_N93_PULSESHAPING_OUT), .A1 (XNOR_1_4_N93_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_6_N93_PULSESHAPING (.ZN (XNOR_1_6_N93_PULSESHAPING_OUT), .A1 (XNOR_1_5_N93_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_7_N93_PULSESHAPING (.ZN (N93), .A1 (XNOR_1_6_N93_PULSESHAPING_OUT), .A2 (GND));

      wire XNOR_1_1_N97_PULSESHAPING_OUT, XNOR_1_2_N97_PULSESHAPING_OUT, XNOR_1_3_N97_PULSESHAPING_OUT, XNOR_1_4_N97_PULSESHAPING_OUT, XNOR_1_5_N97_PULSESHAPING_OUT, XNOR_1_6_N97_PULSESHAPING_OUT;
      NOR2_X1 XNOR_1_1_N97_PULSESHAPING (.ZN (XNOR_1_1_N97_PULSESHAPING_OUT), .A1 (N97_PWL), .A2 (GND));
      NOR2_X1 XNOR_1_2_N97_PULSESHAPING (.ZN (XNOR_1_2_N97_PULSESHAPING_OUT), .A1 (XNOR_1_1_N97_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_3_N97_PULSESHAPING (.ZN (XNOR_1_3_N97_PULSESHAPING_OUT), .A1 (XNOR_1_2_N97_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_4_N97_PULSESHAPING (.ZN (XNOR_1_4_N97_PULSESHAPING_OUT), .A1 (XNOR_1_3_N97_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_5_N97_PULSESHAPING (.ZN (XNOR_1_5_N97_PULSESHAPING_OUT), .A1 (XNOR_1_4_N97_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_6_N97_PULSESHAPING (.ZN (XNOR_1_6_N97_PULSESHAPING_OUT), .A1 (XNOR_1_5_N97_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_7_N97_PULSESHAPING (.ZN (N97), .A1 (XNOR_1_6_N97_PULSESHAPING_OUT), .A2 (GND));

      wire XNOR_1_1_N101_PULSESHAPING_OUT, XNOR_1_2_N101_PULSESHAPING_OUT, XNOR_1_3_N101_PULSESHAPING_OUT, XNOR_1_4_N101_PULSESHAPING_OUT, XNOR_1_5_N101_PULSESHAPING_OUT, XNOR_1_6_N101_PULSESHAPING_OUT;
      NOR2_X1 XNOR_1_1_N101_PULSESHAPING (.ZN (XNOR_1_1_N101_PULSESHAPING_OUT), .A1 (N101_PWL), .A2 (GND));
      NOR2_X1 XNOR_1_2_N101_PULSESHAPING (.ZN (XNOR_1_2_N101_PULSESHAPING_OUT), .A1 (XNOR_1_1_N101_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_3_N101_PULSESHAPING (.ZN (XNOR_1_3_N101_PULSESHAPING_OUT), .A1 (XNOR_1_2_N101_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_4_N101_PULSESHAPING (.ZN (XNOR_1_4_N101_PULSESHAPING_OUT), .A1 (XNOR_1_3_N101_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_5_N101_PULSESHAPING (.ZN (XNOR_1_5_N101_PULSESHAPING_OUT), .A1 (XNOR_1_4_N101_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_6_N101_PULSESHAPING (.ZN (XNOR_1_6_N101_PULSESHAPING_OUT), .A1 (XNOR_1_5_N101_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_7_N101_PULSESHAPING (.ZN (N101), .A1 (XNOR_1_6_N101_PULSESHAPING_OUT), .A2 (GND));

      wire XNOR_1_1_N105_PULSESHAPING_OUT, XNOR_1_2_N105_PULSESHAPING_OUT, XNOR_1_3_N105_PULSESHAPING_OUT, XNOR_1_4_N105_PULSESHAPING_OUT, XNOR_1_5_N105_PULSESHAPING_OUT, XNOR_1_6_N105_PULSESHAPING_OUT;
      NOR2_X1 XNOR_1_1_N105_PULSESHAPING (.ZN (XNOR_1_1_N105_PULSESHAPING_OUT), .A1 (N105_PWL), .A2 (GND));
      NOR2_X1 XNOR_1_2_N105_PULSESHAPING (.ZN (XNOR_1_2_N105_PULSESHAPING_OUT), .A1 (XNOR_1_1_N105_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_3_N105_PULSESHAPING (.ZN (XNOR_1_3_N105_PULSESHAPING_OUT), .A1 (XNOR_1_2_N105_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_4_N105_PULSESHAPING (.ZN (XNOR_1_4_N105_PULSESHAPING_OUT), .A1 (XNOR_1_3_N105_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_5_N105_PULSESHAPING (.ZN (XNOR_1_5_N105_PULSESHAPING_OUT), .A1 (XNOR_1_4_N105_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_6_N105_PULSESHAPING (.ZN (XNOR_1_6_N105_PULSESHAPING_OUT), .A1 (XNOR_1_5_N105_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_7_N105_PULSESHAPING (.ZN (N105), .A1 (XNOR_1_6_N105_PULSESHAPING_OUT), .A2 (GND));

      wire XNOR_1_1_N109_PULSESHAPING_OUT, XNOR_1_2_N109_PULSESHAPING_OUT, XNOR_1_3_N109_PULSESHAPING_OUT, XNOR_1_4_N109_PULSESHAPING_OUT, XNOR_1_5_N109_PULSESHAPING_OUT, XNOR_1_6_N109_PULSESHAPING_OUT;
      NOR2_X1 XNOR_1_1_N109_PULSESHAPING (.ZN (XNOR_1_1_N109_PULSESHAPING_OUT), .A1 (N109_PWL), .A2 (GND));
      NOR2_X1 XNOR_1_2_N109_PULSESHAPING (.ZN (XNOR_1_2_N109_PULSESHAPING_OUT), .A1 (XNOR_1_1_N109_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_3_N109_PULSESHAPING (.ZN (XNOR_1_3_N109_PULSESHAPING_OUT), .A1 (XNOR_1_2_N109_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_4_N109_PULSESHAPING (.ZN (XNOR_1_4_N109_PULSESHAPING_OUT), .A1 (XNOR_1_3_N109_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_5_N109_PULSESHAPING (.ZN (XNOR_1_5_N109_PULSESHAPING_OUT), .A1 (XNOR_1_4_N109_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_6_N109_PULSESHAPING (.ZN (XNOR_1_6_N109_PULSESHAPING_OUT), .A1 (XNOR_1_5_N109_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_7_N109_PULSESHAPING (.ZN (N109), .A1 (XNOR_1_6_N109_PULSESHAPING_OUT), .A2 (GND));

      wire XNOR_1_1_N113_PULSESHAPING_OUT, XNOR_1_2_N113_PULSESHAPING_OUT, XNOR_1_3_N113_PULSESHAPING_OUT, XNOR_1_4_N113_PULSESHAPING_OUT, XNOR_1_5_N113_PULSESHAPING_OUT, XNOR_1_6_N113_PULSESHAPING_OUT;
      NOR2_X1 XNOR_1_1_N113_PULSESHAPING (.ZN (XNOR_1_1_N113_PULSESHAPING_OUT), .A1 (N113_PWL), .A2 (GND));
      NOR2_X1 XNOR_1_2_N113_PULSESHAPING (.ZN (XNOR_1_2_N113_PULSESHAPING_OUT), .A1 (XNOR_1_1_N113_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_3_N113_PULSESHAPING (.ZN (XNOR_1_3_N113_PULSESHAPING_OUT), .A1 (XNOR_1_2_N113_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_4_N113_PULSESHAPING (.ZN (XNOR_1_4_N113_PULSESHAPING_OUT), .A1 (XNOR_1_3_N113_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_5_N113_PULSESHAPING (.ZN (XNOR_1_5_N113_PULSESHAPING_OUT), .A1 (XNOR_1_4_N113_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_6_N113_PULSESHAPING (.ZN (XNOR_1_6_N113_PULSESHAPING_OUT), .A1 (XNOR_1_5_N113_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_7_N113_PULSESHAPING (.ZN (N113), .A1 (XNOR_1_6_N113_PULSESHAPING_OUT), .A2 (GND));

      wire XNOR_1_1_N117_PULSESHAPING_OUT, XNOR_1_2_N117_PULSESHAPING_OUT, XNOR_1_3_N117_PULSESHAPING_OUT, XNOR_1_4_N117_PULSESHAPING_OUT, XNOR_1_5_N117_PULSESHAPING_OUT, XNOR_1_6_N117_PULSESHAPING_OUT;
      NOR2_X1 XNOR_1_1_N117_PULSESHAPING (.ZN (XNOR_1_1_N117_PULSESHAPING_OUT), .A1 (N117_PWL), .A2 (GND));
      NOR2_X1 XNOR_1_2_N117_PULSESHAPING (.ZN (XNOR_1_2_N117_PULSESHAPING_OUT), .A1 (XNOR_1_1_N117_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_3_N117_PULSESHAPING (.ZN (XNOR_1_3_N117_PULSESHAPING_OUT), .A1 (XNOR_1_2_N117_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_4_N117_PULSESHAPING (.ZN (XNOR_1_4_N117_PULSESHAPING_OUT), .A1 (XNOR_1_3_N117_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_5_N117_PULSESHAPING (.ZN (XNOR_1_5_N117_PULSESHAPING_OUT), .A1 (XNOR_1_4_N117_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_6_N117_PULSESHAPING (.ZN (XNOR_1_6_N117_PULSESHAPING_OUT), .A1 (XNOR_1_5_N117_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_7_N117_PULSESHAPING (.ZN (N117), .A1 (XNOR_1_6_N117_PULSESHAPING_OUT), .A2 (GND));

      wire XNOR_1_1_N121_PULSESHAPING_OUT, XNOR_1_2_N121_PULSESHAPING_OUT, XNOR_1_3_N121_PULSESHAPING_OUT, XNOR_1_4_N121_PULSESHAPING_OUT, XNOR_1_5_N121_PULSESHAPING_OUT, XNOR_1_6_N121_PULSESHAPING_OUT;
      NOR2_X1 XNOR_1_1_N121_PULSESHAPING (.ZN (XNOR_1_1_N121_PULSESHAPING_OUT), .A1 (N121_PWL), .A2 (GND));
      NOR2_X1 XNOR_1_2_N121_PULSESHAPING (.ZN (XNOR_1_2_N121_PULSESHAPING_OUT), .A1 (XNOR_1_1_N121_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_3_N121_PULSESHAPING (.ZN (XNOR_1_3_N121_PULSESHAPING_OUT), .A1 (XNOR_1_2_N121_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_4_N121_PULSESHAPING (.ZN (XNOR_1_4_N121_PULSESHAPING_OUT), .A1 (XNOR_1_3_N121_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_5_N121_PULSESHAPING (.ZN (XNOR_1_5_N121_PULSESHAPING_OUT), .A1 (XNOR_1_4_N121_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_6_N121_PULSESHAPING (.ZN (XNOR_1_6_N121_PULSESHAPING_OUT), .A1 (XNOR_1_5_N121_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_7_N121_PULSESHAPING (.ZN (N121), .A1 (XNOR_1_6_N121_PULSESHAPING_OUT), .A2 (GND));

      wire XNOR_1_1_N125_PULSESHAPING_OUT, XNOR_1_2_N125_PULSESHAPING_OUT, XNOR_1_3_N125_PULSESHAPING_OUT, XNOR_1_4_N125_PULSESHAPING_OUT, XNOR_1_5_N125_PULSESHAPING_OUT, XNOR_1_6_N125_PULSESHAPING_OUT;
      NOR2_X1 XNOR_1_1_N125_PULSESHAPING (.ZN (XNOR_1_1_N125_PULSESHAPING_OUT), .A1 (N125_PWL), .A2 (GND));
      NOR2_X1 XNOR_1_2_N125_PULSESHAPING (.ZN (XNOR_1_2_N125_PULSESHAPING_OUT), .A1 (XNOR_1_1_N125_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_3_N125_PULSESHAPING (.ZN (XNOR_1_3_N125_PULSESHAPING_OUT), .A1 (XNOR_1_2_N125_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_4_N125_PULSESHAPING (.ZN (XNOR_1_4_N125_PULSESHAPING_OUT), .A1 (XNOR_1_3_N125_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_5_N125_PULSESHAPING (.ZN (XNOR_1_5_N125_PULSESHAPING_OUT), .A1 (XNOR_1_4_N125_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_6_N125_PULSESHAPING (.ZN (XNOR_1_6_N125_PULSESHAPING_OUT), .A1 (XNOR_1_5_N125_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_7_N125_PULSESHAPING (.ZN (N125), .A1 (XNOR_1_6_N125_PULSESHAPING_OUT), .A2 (GND));

      wire XNOR_1_1_N129_PULSESHAPING_OUT, XNOR_1_2_N129_PULSESHAPING_OUT, XNOR_1_3_N129_PULSESHAPING_OUT, XNOR_1_4_N129_PULSESHAPING_OUT, XNOR_1_5_N129_PULSESHAPING_OUT, XNOR_1_6_N129_PULSESHAPING_OUT;
      NOR2_X1 XNOR_1_1_N129_PULSESHAPING (.ZN (XNOR_1_1_N129_PULSESHAPING_OUT), .A1 (N129_PWL), .A2 (GND));
      NOR2_X1 XNOR_1_2_N129_PULSESHAPING (.ZN (XNOR_1_2_N129_PULSESHAPING_OUT), .A1 (XNOR_1_1_N129_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_3_N129_PULSESHAPING (.ZN (XNOR_1_3_N129_PULSESHAPING_OUT), .A1 (XNOR_1_2_N129_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_4_N129_PULSESHAPING (.ZN (XNOR_1_4_N129_PULSESHAPING_OUT), .A1 (XNOR_1_3_N129_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_5_N129_PULSESHAPING (.ZN (XNOR_1_5_N129_PULSESHAPING_OUT), .A1 (XNOR_1_4_N129_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_6_N129_PULSESHAPING (.ZN (XNOR_1_6_N129_PULSESHAPING_OUT), .A1 (XNOR_1_5_N129_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_7_N129_PULSESHAPING (.ZN (N129), .A1 (XNOR_1_6_N129_PULSESHAPING_OUT), .A2 (GND));

      wire XNOR_1_1_N130_PULSESHAPING_OUT, XNOR_1_2_N130_PULSESHAPING_OUT, XNOR_1_3_N130_PULSESHAPING_OUT, XNOR_1_4_N130_PULSESHAPING_OUT, XNOR_1_5_N130_PULSESHAPING_OUT, XNOR_1_6_N130_PULSESHAPING_OUT;
      NOR2_X1 XNOR_1_1_N130_PULSESHAPING (.ZN (XNOR_1_1_N130_PULSESHAPING_OUT), .A1 (N130_PWL), .A2 (GND));
      NOR2_X1 XNOR_1_2_N130_PULSESHAPING (.ZN (XNOR_1_2_N130_PULSESHAPING_OUT), .A1 (XNOR_1_1_N130_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_3_N130_PULSESHAPING (.ZN (XNOR_1_3_N130_PULSESHAPING_OUT), .A1 (XNOR_1_2_N130_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_4_N130_PULSESHAPING (.ZN (XNOR_1_4_N130_PULSESHAPING_OUT), .A1 (XNOR_1_3_N130_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_5_N130_PULSESHAPING (.ZN (XNOR_1_5_N130_PULSESHAPING_OUT), .A1 (XNOR_1_4_N130_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_6_N130_PULSESHAPING (.ZN (XNOR_1_6_N130_PULSESHAPING_OUT), .A1 (XNOR_1_5_N130_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_7_N130_PULSESHAPING (.ZN (N130), .A1 (XNOR_1_6_N130_PULSESHAPING_OUT), .A2 (GND));

      wire XNOR_1_1_N131_PULSESHAPING_OUT, XNOR_1_2_N131_PULSESHAPING_OUT, XNOR_1_3_N131_PULSESHAPING_OUT, XNOR_1_4_N131_PULSESHAPING_OUT, XNOR_1_5_N131_PULSESHAPING_OUT, XNOR_1_6_N131_PULSESHAPING_OUT;
      NOR2_X1 XNOR_1_1_N131_PULSESHAPING (.ZN (XNOR_1_1_N131_PULSESHAPING_OUT), .A1 (N131_PWL), .A2 (GND));
      NOR2_X1 XNOR_1_2_N131_PULSESHAPING (.ZN (XNOR_1_2_N131_PULSESHAPING_OUT), .A1 (XNOR_1_1_N131_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_3_N131_PULSESHAPING (.ZN (XNOR_1_3_N131_PULSESHAPING_OUT), .A1 (XNOR_1_2_N131_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_4_N131_PULSESHAPING (.ZN (XNOR_1_4_N131_PULSESHAPING_OUT), .A1 (XNOR_1_3_N131_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_5_N131_PULSESHAPING (.ZN (XNOR_1_5_N131_PULSESHAPING_OUT), .A1 (XNOR_1_4_N131_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_6_N131_PULSESHAPING (.ZN (XNOR_1_6_N131_PULSESHAPING_OUT), .A1 (XNOR_1_5_N131_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_7_N131_PULSESHAPING (.ZN (N131), .A1 (XNOR_1_6_N131_PULSESHAPING_OUT), .A2 (GND));

      wire XNOR_1_1_N132_PULSESHAPING_OUT, XNOR_1_2_N132_PULSESHAPING_OUT, XNOR_1_3_N132_PULSESHAPING_OUT, XNOR_1_4_N132_PULSESHAPING_OUT, XNOR_1_5_N132_PULSESHAPING_OUT, XNOR_1_6_N132_PULSESHAPING_OUT;
      NOR2_X1 XNOR_1_1_N132_PULSESHAPING (.ZN (XNOR_1_1_N132_PULSESHAPING_OUT), .A1 (N132_PWL), .A2 (GND));
      NOR2_X1 XNOR_1_2_N132_PULSESHAPING (.ZN (XNOR_1_2_N132_PULSESHAPING_OUT), .A1 (XNOR_1_1_N132_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_3_N132_PULSESHAPING (.ZN (XNOR_1_3_N132_PULSESHAPING_OUT), .A1 (XNOR_1_2_N132_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_4_N132_PULSESHAPING (.ZN (XNOR_1_4_N132_PULSESHAPING_OUT), .A1 (XNOR_1_3_N132_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_5_N132_PULSESHAPING (.ZN (XNOR_1_5_N132_PULSESHAPING_OUT), .A1 (XNOR_1_4_N132_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_6_N132_PULSESHAPING (.ZN (XNOR_1_6_N132_PULSESHAPING_OUT), .A1 (XNOR_1_5_N132_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_7_N132_PULSESHAPING (.ZN (N132), .A1 (XNOR_1_6_N132_PULSESHAPING_OUT), .A2 (GND));

      wire XNOR_1_1_N133_PULSESHAPING_OUT, XNOR_1_2_N133_PULSESHAPING_OUT, XNOR_1_3_N133_PULSESHAPING_OUT, XNOR_1_4_N133_PULSESHAPING_OUT, XNOR_1_5_N133_PULSESHAPING_OUT, XNOR_1_6_N133_PULSESHAPING_OUT;
      NOR2_X1 XNOR_1_1_N133_PULSESHAPING (.ZN (XNOR_1_1_N133_PULSESHAPING_OUT), .A1 (N133_PWL), .A2 (GND));
      NOR2_X1 XNOR_1_2_N133_PULSESHAPING (.ZN (XNOR_1_2_N133_PULSESHAPING_OUT), .A1 (XNOR_1_1_N133_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_3_N133_PULSESHAPING (.ZN (XNOR_1_3_N133_PULSESHAPING_OUT), .A1 (XNOR_1_2_N133_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_4_N133_PULSESHAPING (.ZN (XNOR_1_4_N133_PULSESHAPING_OUT), .A1 (XNOR_1_3_N133_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_5_N133_PULSESHAPING (.ZN (XNOR_1_5_N133_PULSESHAPING_OUT), .A1 (XNOR_1_4_N133_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_6_N133_PULSESHAPING (.ZN (XNOR_1_6_N133_PULSESHAPING_OUT), .A1 (XNOR_1_5_N133_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_7_N133_PULSESHAPING (.ZN (N133), .A1 (XNOR_1_6_N133_PULSESHAPING_OUT), .A2 (GND));

      wire XNOR_1_1_N134_PULSESHAPING_OUT, XNOR_1_2_N134_PULSESHAPING_OUT, XNOR_1_3_N134_PULSESHAPING_OUT, XNOR_1_4_N134_PULSESHAPING_OUT, XNOR_1_5_N134_PULSESHAPING_OUT, XNOR_1_6_N134_PULSESHAPING_OUT;
      NOR2_X1 XNOR_1_1_N134_PULSESHAPING (.ZN (XNOR_1_1_N134_PULSESHAPING_OUT), .A1 (N134_PWL), .A2 (GND));
      NOR2_X1 XNOR_1_2_N134_PULSESHAPING (.ZN (XNOR_1_2_N134_PULSESHAPING_OUT), .A1 (XNOR_1_1_N134_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_3_N134_PULSESHAPING (.ZN (XNOR_1_3_N134_PULSESHAPING_OUT), .A1 (XNOR_1_2_N134_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_4_N134_PULSESHAPING (.ZN (XNOR_1_4_N134_PULSESHAPING_OUT), .A1 (XNOR_1_3_N134_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_5_N134_PULSESHAPING (.ZN (XNOR_1_5_N134_PULSESHAPING_OUT), .A1 (XNOR_1_4_N134_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_6_N134_PULSESHAPING (.ZN (XNOR_1_6_N134_PULSESHAPING_OUT), .A1 (XNOR_1_5_N134_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_7_N134_PULSESHAPING (.ZN (N134), .A1 (XNOR_1_6_N134_PULSESHAPING_OUT), .A2 (GND));

      wire XNOR_1_1_N135_PULSESHAPING_OUT, XNOR_1_2_N135_PULSESHAPING_OUT, XNOR_1_3_N135_PULSESHAPING_OUT, XNOR_1_4_N135_PULSESHAPING_OUT, XNOR_1_5_N135_PULSESHAPING_OUT, XNOR_1_6_N135_PULSESHAPING_OUT;
      NOR2_X1 XNOR_1_1_N135_PULSESHAPING (.ZN (XNOR_1_1_N135_PULSESHAPING_OUT), .A1 (N135_PWL), .A2 (GND));
      NOR2_X1 XNOR_1_2_N135_PULSESHAPING (.ZN (XNOR_1_2_N135_PULSESHAPING_OUT), .A1 (XNOR_1_1_N135_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_3_N135_PULSESHAPING (.ZN (XNOR_1_3_N135_PULSESHAPING_OUT), .A1 (XNOR_1_2_N135_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_4_N135_PULSESHAPING (.ZN (XNOR_1_4_N135_PULSESHAPING_OUT), .A1 (XNOR_1_3_N135_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_5_N135_PULSESHAPING (.ZN (XNOR_1_5_N135_PULSESHAPING_OUT), .A1 (XNOR_1_4_N135_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_6_N135_PULSESHAPING (.ZN (XNOR_1_6_N135_PULSESHAPING_OUT), .A1 (XNOR_1_5_N135_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_7_N135_PULSESHAPING (.ZN (N135), .A1 (XNOR_1_6_N135_PULSESHAPING_OUT), .A2 (GND));

      wire XNOR_1_1_N136_PULSESHAPING_OUT, XNOR_1_2_N136_PULSESHAPING_OUT, XNOR_1_3_N136_PULSESHAPING_OUT, XNOR_1_4_N136_PULSESHAPING_OUT, XNOR_1_5_N136_PULSESHAPING_OUT, XNOR_1_6_N136_PULSESHAPING_OUT;
      NOR2_X1 XNOR_1_1_N136_PULSESHAPING (.ZN (XNOR_1_1_N136_PULSESHAPING_OUT), .A1 (N136_PWL), .A2 (GND));
      NOR2_X1 XNOR_1_2_N136_PULSESHAPING (.ZN (XNOR_1_2_N136_PULSESHAPING_OUT), .A1 (XNOR_1_1_N136_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_3_N136_PULSESHAPING (.ZN (XNOR_1_3_N136_PULSESHAPING_OUT), .A1 (XNOR_1_2_N136_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_4_N136_PULSESHAPING (.ZN (XNOR_1_4_N136_PULSESHAPING_OUT), .A1 (XNOR_1_3_N136_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_5_N136_PULSESHAPING (.ZN (XNOR_1_5_N136_PULSESHAPING_OUT), .A1 (XNOR_1_4_N136_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_6_N136_PULSESHAPING (.ZN (XNOR_1_6_N136_PULSESHAPING_OUT), .A1 (XNOR_1_5_N136_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_7_N136_PULSESHAPING (.ZN (N136), .A1 (XNOR_1_6_N136_PULSESHAPING_OUT), .A2 (GND));

      wire XNOR_1_1_N137_PULSESHAPING_OUT, XNOR_1_2_N137_PULSESHAPING_OUT, XNOR_1_3_N137_PULSESHAPING_OUT, XNOR_1_4_N137_PULSESHAPING_OUT, XNOR_1_5_N137_PULSESHAPING_OUT, XNOR_1_6_N137_PULSESHAPING_OUT;
      NOR2_X1 XNOR_1_1_N137_PULSESHAPING (.ZN (XNOR_1_1_N137_PULSESHAPING_OUT), .A1 (N137_PWL), .A2 (GND));
      NOR2_X1 XNOR_1_2_N137_PULSESHAPING (.ZN (XNOR_1_2_N137_PULSESHAPING_OUT), .A1 (XNOR_1_1_N137_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_3_N137_PULSESHAPING (.ZN (XNOR_1_3_N137_PULSESHAPING_OUT), .A1 (XNOR_1_2_N137_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_4_N137_PULSESHAPING (.ZN (XNOR_1_4_N137_PULSESHAPING_OUT), .A1 (XNOR_1_3_N137_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_5_N137_PULSESHAPING (.ZN (XNOR_1_5_N137_PULSESHAPING_OUT), .A1 (XNOR_1_4_N137_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_6_N137_PULSESHAPING (.ZN (XNOR_1_6_N137_PULSESHAPING_OUT), .A1 (XNOR_1_5_N137_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_7_N137_PULSESHAPING (.ZN (N137), .A1 (XNOR_1_6_N137_PULSESHAPING_OUT), .A2 (GND));



      wire XNOR_1_1_NUM1_OUT, XNOR_1_2_NUM1_OUT, XNOR_1_3_NUM1_OUT, XNOR_1_4_NUM1_OUT;
      NOR2_X1 XNOR_1_1_NUM1 (.ZN (XNOR_1_1_NUM1_OUT), .A1 (N1), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM1 (.ZN (XNOR_1_2_NUM1_OUT), .A1 (GND), .A2 (N5));
      NOR2_X1 XNOR_1_3_NUM1 (.ZN (XNOR_1_3_NUM1_OUT), .A1 (XNOR_1_1_NUM1_OUT), .A2 (XNOR_1_2_NUM1_OUT));
      NOR2_X1 XNOR_1_4_NUM1 (.ZN (XNOR_1_4_NUM1_OUT), .A1 (N1), .A2 (N5));
      NOR2_X1 XNOR_1_5_NUM1 (.ZN (N250), .A1 (XNOR_1_3_NUM1_OUT), .A2 (XNOR_1_4_NUM1_OUT));
      wire XNOR_1_1_NUM2_OUT, XNOR_1_2_NUM2_OUT, XNOR_1_3_NUM2_OUT, XNOR_1_4_NUM2_OUT;
      NOR2_X1 XNOR_1_1_NUM2 (.ZN (XNOR_1_1_NUM2_OUT), .A1 (N9), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM2 (.ZN (XNOR_1_2_NUM2_OUT), .A1 (GND), .A2 (N13));
      NOR2_X1 XNOR_1_3_NUM2 (.ZN (XNOR_1_3_NUM2_OUT), .A1 (XNOR_1_1_NUM2_OUT), .A2 (XNOR_1_2_NUM2_OUT));
      NOR2_X1 XNOR_1_4_NUM2 (.ZN (XNOR_1_4_NUM2_OUT), .A1 (N9), .A2 (N13));
      NOR2_X1 XNOR_1_5_NUM2 (.ZN (N251), .A1 (XNOR_1_3_NUM2_OUT), .A2 (XNOR_1_4_NUM2_OUT));
      wire XNOR_1_1_NUM3_OUT, XNOR_1_2_NUM3_OUT, XNOR_1_3_NUM3_OUT, XNOR_1_4_NUM3_OUT;
      NOR2_X1 XNOR_1_1_NUM3 (.ZN (XNOR_1_1_NUM3_OUT), .A1 (N17), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM3 (.ZN (XNOR_1_2_NUM3_OUT), .A1 (GND), .A2 (N21));
      NOR2_X1 XNOR_1_3_NUM3 (.ZN (XNOR_1_3_NUM3_OUT), .A1 (XNOR_1_1_NUM3_OUT), .A2 (XNOR_1_2_NUM3_OUT));
      NOR2_X1 XNOR_1_4_NUM3 (.ZN (XNOR_1_4_NUM3_OUT), .A1 (N17), .A2 (N21));
      NOR2_X1 XNOR_1_5_NUM3 (.ZN (N252), .A1 (XNOR_1_3_NUM3_OUT), .A2 (XNOR_1_4_NUM3_OUT));
      wire XNOR_1_1_NUM4_OUT, XNOR_1_2_NUM4_OUT, XNOR_1_3_NUM4_OUT, XNOR_1_4_NUM4_OUT;
      NOR2_X1 XNOR_1_1_NUM4 (.ZN (XNOR_1_1_NUM4_OUT), .A1 (N25), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM4 (.ZN (XNOR_1_2_NUM4_OUT), .A1 (GND), .A2 (N29));
      NOR2_X1 XNOR_1_3_NUM4 (.ZN (XNOR_1_3_NUM4_OUT), .A1 (XNOR_1_1_NUM4_OUT), .A2 (XNOR_1_2_NUM4_OUT));
      NOR2_X1 XNOR_1_4_NUM4 (.ZN (XNOR_1_4_NUM4_OUT), .A1 (N25), .A2 (N29));
      NOR2_X1 XNOR_1_5_NUM4 (.ZN (N253), .A1 (XNOR_1_3_NUM4_OUT), .A2 (XNOR_1_4_NUM4_OUT));
      wire XNOR_1_1_NUM5_OUT, XNOR_1_2_NUM5_OUT, XNOR_1_3_NUM5_OUT, XNOR_1_4_NUM5_OUT;
      NOR2_X1 XNOR_1_1_NUM5 (.ZN (XNOR_1_1_NUM5_OUT), .A1 (N33), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM5 (.ZN (XNOR_1_2_NUM5_OUT), .A1 (GND), .A2 (N37));
      NOR2_X1 XNOR_1_3_NUM5 (.ZN (XNOR_1_3_NUM5_OUT), .A1 (XNOR_1_1_NUM5_OUT), .A2 (XNOR_1_2_NUM5_OUT));
      NOR2_X1 XNOR_1_4_NUM5 (.ZN (XNOR_1_4_NUM5_OUT), .A1 (N33), .A2 (N37));
      NOR2_X1 XNOR_1_5_NUM5 (.ZN (N254), .A1 (XNOR_1_3_NUM5_OUT), .A2 (XNOR_1_4_NUM5_OUT));
      wire XNOR_1_1_NUM6_OUT, XNOR_1_2_NUM6_OUT, XNOR_1_3_NUM6_OUT, XNOR_1_4_NUM6_OUT;
      NOR2_X1 XNOR_1_1_NUM6 (.ZN (XNOR_1_1_NUM6_OUT), .A1 (N41), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM6 (.ZN (XNOR_1_2_NUM6_OUT), .A1 (GND), .A2 (N45));
      NOR2_X1 XNOR_1_3_NUM6 (.ZN (XNOR_1_3_NUM6_OUT), .A1 (XNOR_1_1_NUM6_OUT), .A2 (XNOR_1_2_NUM6_OUT));
      NOR2_X1 XNOR_1_4_NUM6 (.ZN (XNOR_1_4_NUM6_OUT), .A1 (N41), .A2 (N45));
      NOR2_X1 XNOR_1_5_NUM6 (.ZN (N255), .A1 (XNOR_1_3_NUM6_OUT), .A2 (XNOR_1_4_NUM6_OUT));
      wire XNOR_1_1_NUM7_OUT, XNOR_1_2_NUM7_OUT, XNOR_1_3_NUM7_OUT, XNOR_1_4_NUM7_OUT;
      NOR2_X1 XNOR_1_1_NUM7 (.ZN (XNOR_1_1_NUM7_OUT), .A1 (N49), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM7 (.ZN (XNOR_1_2_NUM7_OUT), .A1 (GND), .A2 (N53));
      NOR2_X1 XNOR_1_3_NUM7 (.ZN (XNOR_1_3_NUM7_OUT), .A1 (XNOR_1_1_NUM7_OUT), .A2 (XNOR_1_2_NUM7_OUT));
      NOR2_X1 XNOR_1_4_NUM7 (.ZN (XNOR_1_4_NUM7_OUT), .A1 (N49), .A2 (N53));
      NOR2_X1 XNOR_1_5_NUM7 (.ZN (N256), .A1 (XNOR_1_3_NUM7_OUT), .A2 (XNOR_1_4_NUM7_OUT));
      wire XNOR_1_1_NUM8_OUT, XNOR_1_2_NUM8_OUT, XNOR_1_3_NUM8_OUT, XNOR_1_4_NUM8_OUT;
      NOR2_X1 XNOR_1_1_NUM8 (.ZN (XNOR_1_1_NUM8_OUT), .A1 (N57), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM8 (.ZN (XNOR_1_2_NUM8_OUT), .A1 (GND), .A2 (N61));
      NOR2_X1 XNOR_1_3_NUM8 (.ZN (XNOR_1_3_NUM8_OUT), .A1 (XNOR_1_1_NUM8_OUT), .A2 (XNOR_1_2_NUM8_OUT));
      NOR2_X1 XNOR_1_4_NUM8 (.ZN (XNOR_1_4_NUM8_OUT), .A1 (N57), .A2 (N61));
      NOR2_X1 XNOR_1_5_NUM8 (.ZN (N257), .A1 (XNOR_1_3_NUM8_OUT), .A2 (XNOR_1_4_NUM8_OUT));
      wire XNOR_1_1_NUM9_OUT, XNOR_1_2_NUM9_OUT, XNOR_1_3_NUM9_OUT, XNOR_1_4_NUM9_OUT;
      NOR2_X1 XNOR_1_1_NUM9 (.ZN (XNOR_1_1_NUM9_OUT), .A1 (N65), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM9 (.ZN (XNOR_1_2_NUM9_OUT), .A1 (GND), .A2 (N69));
      NOR2_X1 XNOR_1_3_NUM9 (.ZN (XNOR_1_3_NUM9_OUT), .A1 (XNOR_1_1_NUM9_OUT), .A2 (XNOR_1_2_NUM9_OUT));
      NOR2_X1 XNOR_1_4_NUM9 (.ZN (XNOR_1_4_NUM9_OUT), .A1 (N65), .A2 (N69));
      NOR2_X1 XNOR_1_5_NUM9 (.ZN (N258), .A1 (XNOR_1_3_NUM9_OUT), .A2 (XNOR_1_4_NUM9_OUT));
      wire XNOR_1_1_NUM10_OUT, XNOR_1_2_NUM10_OUT, XNOR_1_3_NUM10_OUT, XNOR_1_4_NUM10_OUT;
      NOR2_X1 XNOR_1_1_NUM10 (.ZN (XNOR_1_1_NUM10_OUT), .A1 (N73), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM10 (.ZN (XNOR_1_2_NUM10_OUT), .A1 (GND), .A2 (N77));
      NOR2_X1 XNOR_1_3_NUM10 (.ZN (XNOR_1_3_NUM10_OUT), .A1 (XNOR_1_1_NUM10_OUT), .A2 (XNOR_1_2_NUM10_OUT));
      NOR2_X1 XNOR_1_4_NUM10 (.ZN (XNOR_1_4_NUM10_OUT), .A1 (N73), .A2 (N77));
      NOR2_X1 XNOR_1_5_NUM10 (.ZN (N259), .A1 (XNOR_1_3_NUM10_OUT), .A2 (XNOR_1_4_NUM10_OUT));
      wire XNOR_1_1_NUM11_OUT, XNOR_1_2_NUM11_OUT, XNOR_1_3_NUM11_OUT, XNOR_1_4_NUM11_OUT;
      NOR2_X1 XNOR_1_1_NUM11 (.ZN (XNOR_1_1_NUM11_OUT), .A1 (N81), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM11 (.ZN (XNOR_1_2_NUM11_OUT), .A1 (GND), .A2 (N85));
      NOR2_X1 XNOR_1_3_NUM11 (.ZN (XNOR_1_3_NUM11_OUT), .A1 (XNOR_1_1_NUM11_OUT), .A2 (XNOR_1_2_NUM11_OUT));
      NOR2_X1 XNOR_1_4_NUM11 (.ZN (XNOR_1_4_NUM11_OUT), .A1 (N81), .A2 (N85));
      NOR2_X1 XNOR_1_5_NUM11 (.ZN (N260), .A1 (XNOR_1_3_NUM11_OUT), .A2 (XNOR_1_4_NUM11_OUT));
      wire XNOR_1_1_NUM12_OUT, XNOR_1_2_NUM12_OUT, XNOR_1_3_NUM12_OUT, XNOR_1_4_NUM12_OUT;
      NOR2_X1 XNOR_1_1_NUM12 (.ZN (XNOR_1_1_NUM12_OUT), .A1 (N89), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM12 (.ZN (XNOR_1_2_NUM12_OUT), .A1 (GND), .A2 (N93));
      NOR2_X1 XNOR_1_3_NUM12 (.ZN (XNOR_1_3_NUM12_OUT), .A1 (XNOR_1_1_NUM12_OUT), .A2 (XNOR_1_2_NUM12_OUT));
      NOR2_X1 XNOR_1_4_NUM12 (.ZN (XNOR_1_4_NUM12_OUT), .A1 (N89), .A2 (N93));
      NOR2_X1 XNOR_1_5_NUM12 (.ZN (N261), .A1 (XNOR_1_3_NUM12_OUT), .A2 (XNOR_1_4_NUM12_OUT));
      wire XNOR_1_1_NUM13_OUT, XNOR_1_2_NUM13_OUT, XNOR_1_3_NUM13_OUT, XNOR_1_4_NUM13_OUT;
      NOR2_X1 XNOR_1_1_NUM13 (.ZN (XNOR_1_1_NUM13_OUT), .A1 (N97), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM13 (.ZN (XNOR_1_2_NUM13_OUT), .A1 (GND), .A2 (N101));
      NOR2_X1 XNOR_1_3_NUM13 (.ZN (XNOR_1_3_NUM13_OUT), .A1 (XNOR_1_1_NUM13_OUT), .A2 (XNOR_1_2_NUM13_OUT));
      NOR2_X1 XNOR_1_4_NUM13 (.ZN (XNOR_1_4_NUM13_OUT), .A1 (N97), .A2 (N101));
      NOR2_X1 XNOR_1_5_NUM13 (.ZN (N262), .A1 (XNOR_1_3_NUM13_OUT), .A2 (XNOR_1_4_NUM13_OUT));
      wire XNOR_1_1_NUM14_OUT, XNOR_1_2_NUM14_OUT, XNOR_1_3_NUM14_OUT, XNOR_1_4_NUM14_OUT;
      NOR2_X1 XNOR_1_1_NUM14 (.ZN (XNOR_1_1_NUM14_OUT), .A1 (N105), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM14 (.ZN (XNOR_1_2_NUM14_OUT), .A1 (GND), .A2 (N109));
      NOR2_X1 XNOR_1_3_NUM14 (.ZN (XNOR_1_3_NUM14_OUT), .A1 (XNOR_1_1_NUM14_OUT), .A2 (XNOR_1_2_NUM14_OUT));
      NOR2_X1 XNOR_1_4_NUM14 (.ZN (XNOR_1_4_NUM14_OUT), .A1 (N105), .A2 (N109));
      NOR2_X1 XNOR_1_5_NUM14 (.ZN (N263), .A1 (XNOR_1_3_NUM14_OUT), .A2 (XNOR_1_4_NUM14_OUT));
      wire XNOR_1_1_NUM15_OUT, XNOR_1_2_NUM15_OUT, XNOR_1_3_NUM15_OUT, XNOR_1_4_NUM15_OUT;
      NOR2_X1 XNOR_1_1_NUM15 (.ZN (XNOR_1_1_NUM15_OUT), .A1 (N113), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM15 (.ZN (XNOR_1_2_NUM15_OUT), .A1 (GND), .A2 (N117));
      NOR2_X1 XNOR_1_3_NUM15 (.ZN (XNOR_1_3_NUM15_OUT), .A1 (XNOR_1_1_NUM15_OUT), .A2 (XNOR_1_2_NUM15_OUT));
      NOR2_X1 XNOR_1_4_NUM15 (.ZN (XNOR_1_4_NUM15_OUT), .A1 (N113), .A2 (N117));
      NOR2_X1 XNOR_1_5_NUM15 (.ZN (N264), .A1 (XNOR_1_3_NUM15_OUT), .A2 (XNOR_1_4_NUM15_OUT));
      wire XNOR_1_1_NUM16_OUT, XNOR_1_2_NUM16_OUT, XNOR_1_3_NUM16_OUT, XNOR_1_4_NUM16_OUT;
      NOR2_X1 XNOR_1_1_NUM16 (.ZN (XNOR_1_1_NUM16_OUT), .A1 (N121), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM16 (.ZN (XNOR_1_2_NUM16_OUT), .A1 (GND), .A2 (N125));
      NOR2_X1 XNOR_1_3_NUM16 (.ZN (XNOR_1_3_NUM16_OUT), .A1 (XNOR_1_1_NUM16_OUT), .A2 (XNOR_1_2_NUM16_OUT));
      NOR2_X1 XNOR_1_4_NUM16 (.ZN (XNOR_1_4_NUM16_OUT), .A1 (N121), .A2 (N125));
      NOR2_X1 XNOR_1_5_NUM16 (.ZN (N265), .A1 (XNOR_1_3_NUM16_OUT), .A2 (XNOR_1_4_NUM16_OUT));
      wire XNOR_1_1_NUM17_OUT, XNOR_1_2_NUM17_OUT;
      NOR2_X1 XNOR_1_1_NUM17 (.ZN (XNOR_1_1_NUM17_OUT), .A1 (N129), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM17 (.ZN (XNOR_1_2_NUM17_OUT), .A1 (GND), .A2 (N137));
      NOR2_X1 XNOR_1_3_NUM17 (.ZN (N266), .A1 (XNOR_1_1_NUM17_OUT), .A2 (XNOR_1_2_NUM17_OUT));
      wire XNOR_1_1_NUM18_OUT, XNOR_1_2_NUM18_OUT;
      NOR2_X1 XNOR_1_1_NUM18 (.ZN (XNOR_1_1_NUM18_OUT), .A1 (N130), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM18 (.ZN (XNOR_1_2_NUM18_OUT), .A1 (GND), .A2 (N137));
      NOR2_X1 XNOR_1_3_NUM18 (.ZN (N267), .A1 (XNOR_1_1_NUM18_OUT), .A2 (XNOR_1_2_NUM18_OUT));
      wire XNOR_1_1_NUM19_OUT, XNOR_1_2_NUM19_OUT;
      NOR2_X1 XNOR_1_1_NUM19 (.ZN (XNOR_1_1_NUM19_OUT), .A1 (N131), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM19 (.ZN (XNOR_1_2_NUM19_OUT), .A1 (GND), .A2 (N137));
      NOR2_X1 XNOR_1_3_NUM19 (.ZN (N268), .A1 (XNOR_1_1_NUM19_OUT), .A2 (XNOR_1_2_NUM19_OUT));
      wire XNOR_1_1_NUM20_OUT, XNOR_1_2_NUM20_OUT;
      NOR2_X1 XNOR_1_1_NUM20 (.ZN (XNOR_1_1_NUM20_OUT), .A1 (N132), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM20 (.ZN (XNOR_1_2_NUM20_OUT), .A1 (GND), .A2 (N137));
      NOR2_X1 XNOR_1_3_NUM20 (.ZN (N269), .A1 (XNOR_1_1_NUM20_OUT), .A2 (XNOR_1_2_NUM20_OUT));
      wire XNOR_1_1_NUM21_OUT, XNOR_1_2_NUM21_OUT;
      NOR2_X1 XNOR_1_1_NUM21 (.ZN (XNOR_1_1_NUM21_OUT), .A1 (N133), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM21 (.ZN (XNOR_1_2_NUM21_OUT), .A1 (GND), .A2 (N137));
      NOR2_X1 XNOR_1_3_NUM21 (.ZN (N270), .A1 (XNOR_1_1_NUM21_OUT), .A2 (XNOR_1_2_NUM21_OUT));
      wire XNOR_1_1_NUM22_OUT, XNOR_1_2_NUM22_OUT;
      NOR2_X1 XNOR_1_1_NUM22 (.ZN (XNOR_1_1_NUM22_OUT), .A1 (N134), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM22 (.ZN (XNOR_1_2_NUM22_OUT), .A1 (GND), .A2 (N137));
      NOR2_X1 XNOR_1_3_NUM22 (.ZN (N271), .A1 (XNOR_1_1_NUM22_OUT), .A2 (XNOR_1_2_NUM22_OUT));
      wire XNOR_1_1_NUM23_OUT, XNOR_1_2_NUM23_OUT;
      NOR2_X1 XNOR_1_1_NUM23 (.ZN (XNOR_1_1_NUM23_OUT), .A1 (N135), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM23 (.ZN (XNOR_1_2_NUM23_OUT), .A1 (GND), .A2 (N137));
      NOR2_X1 XNOR_1_3_NUM23 (.ZN (N272), .A1 (XNOR_1_1_NUM23_OUT), .A2 (XNOR_1_2_NUM23_OUT));
      wire XNOR_1_1_NUM24_OUT, XNOR_1_2_NUM24_OUT;
      NOR2_X1 XNOR_1_1_NUM24 (.ZN (XNOR_1_1_NUM24_OUT), .A1 (N136), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM24 (.ZN (XNOR_1_2_NUM24_OUT), .A1 (GND), .A2 (N137));
      NOR2_X1 XNOR_1_3_NUM24 (.ZN (N273), .A1 (XNOR_1_1_NUM24_OUT), .A2 (XNOR_1_2_NUM24_OUT));
      wire XNOR_1_1_NUM25_OUT, XNOR_1_2_NUM25_OUT, XNOR_1_3_NUM25_OUT, XNOR_1_4_NUM25_OUT;
      NOR2_X1 XNOR_1_1_NUM25 (.ZN (XNOR_1_1_NUM25_OUT), .A1 (N1), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM25 (.ZN (XNOR_1_2_NUM25_OUT), .A1 (GND), .A2 (N17));
      NOR2_X1 XNOR_1_3_NUM25 (.ZN (XNOR_1_3_NUM25_OUT), .A1 (XNOR_1_1_NUM25_OUT), .A2 (XNOR_1_2_NUM25_OUT));
      NOR2_X1 XNOR_1_4_NUM25 (.ZN (XNOR_1_4_NUM25_OUT), .A1 (N1), .A2 (N17));
      NOR2_X1 XNOR_1_5_NUM25 (.ZN (N274), .A1 (XNOR_1_3_NUM25_OUT), .A2 (XNOR_1_4_NUM25_OUT));
      wire XNOR_1_1_NUM26_OUT, XNOR_1_2_NUM26_OUT, XNOR_1_3_NUM26_OUT, XNOR_1_4_NUM26_OUT;
      NOR2_X1 XNOR_1_1_NUM26 (.ZN (XNOR_1_1_NUM26_OUT), .A1 (N33), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM26 (.ZN (XNOR_1_2_NUM26_OUT), .A1 (GND), .A2 (N49));
      NOR2_X1 XNOR_1_3_NUM26 (.ZN (XNOR_1_3_NUM26_OUT), .A1 (XNOR_1_1_NUM26_OUT), .A2 (XNOR_1_2_NUM26_OUT));
      NOR2_X1 XNOR_1_4_NUM26 (.ZN (XNOR_1_4_NUM26_OUT), .A1 (N33), .A2 (N49));
      NOR2_X1 XNOR_1_5_NUM26 (.ZN (N275), .A1 (XNOR_1_3_NUM26_OUT), .A2 (XNOR_1_4_NUM26_OUT));
      wire XNOR_1_1_NUM27_OUT, XNOR_1_2_NUM27_OUT, XNOR_1_3_NUM27_OUT, XNOR_1_4_NUM27_OUT;
      NOR2_X1 XNOR_1_1_NUM27 (.ZN (XNOR_1_1_NUM27_OUT), .A1 (N5), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM27 (.ZN (XNOR_1_2_NUM27_OUT), .A1 (GND), .A2 (N21));
      NOR2_X1 XNOR_1_3_NUM27 (.ZN (XNOR_1_3_NUM27_OUT), .A1 (XNOR_1_1_NUM27_OUT), .A2 (XNOR_1_2_NUM27_OUT));
      NOR2_X1 XNOR_1_4_NUM27 (.ZN (XNOR_1_4_NUM27_OUT), .A1 (N5), .A2 (N21));
      NOR2_X1 XNOR_1_5_NUM27 (.ZN (N276), .A1 (XNOR_1_3_NUM27_OUT), .A2 (XNOR_1_4_NUM27_OUT));
      wire XNOR_1_1_NUM28_OUT, XNOR_1_2_NUM28_OUT, XNOR_1_3_NUM28_OUT, XNOR_1_4_NUM28_OUT;
      NOR2_X1 XNOR_1_1_NUM28 (.ZN (XNOR_1_1_NUM28_OUT), .A1 (N37), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM28 (.ZN (XNOR_1_2_NUM28_OUT), .A1 (GND), .A2 (N53));
      NOR2_X1 XNOR_1_3_NUM28 (.ZN (XNOR_1_3_NUM28_OUT), .A1 (XNOR_1_1_NUM28_OUT), .A2 (XNOR_1_2_NUM28_OUT));
      NOR2_X1 XNOR_1_4_NUM28 (.ZN (XNOR_1_4_NUM28_OUT), .A1 (N37), .A2 (N53));
      NOR2_X1 XNOR_1_5_NUM28 (.ZN (N277), .A1 (XNOR_1_3_NUM28_OUT), .A2 (XNOR_1_4_NUM28_OUT));
      wire XNOR_1_1_NUM29_OUT, XNOR_1_2_NUM29_OUT, XNOR_1_3_NUM29_OUT, XNOR_1_4_NUM29_OUT;
      NOR2_X1 XNOR_1_1_NUM29 (.ZN (XNOR_1_1_NUM29_OUT), .A1 (N9), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM29 (.ZN (XNOR_1_2_NUM29_OUT), .A1 (GND), .A2 (N25));
      NOR2_X1 XNOR_1_3_NUM29 (.ZN (XNOR_1_3_NUM29_OUT), .A1 (XNOR_1_1_NUM29_OUT), .A2 (XNOR_1_2_NUM29_OUT));
      NOR2_X1 XNOR_1_4_NUM29 (.ZN (XNOR_1_4_NUM29_OUT), .A1 (N9), .A2 (N25));
      NOR2_X1 XNOR_1_5_NUM29 (.ZN (N278), .A1 (XNOR_1_3_NUM29_OUT), .A2 (XNOR_1_4_NUM29_OUT));
      wire XNOR_1_1_NUM30_OUT, XNOR_1_2_NUM30_OUT, XNOR_1_3_NUM30_OUT, XNOR_1_4_NUM30_OUT;
      NOR2_X1 XNOR_1_1_NUM30 (.ZN (XNOR_1_1_NUM30_OUT), .A1 (N41), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM30 (.ZN (XNOR_1_2_NUM30_OUT), .A1 (GND), .A2 (N57));
      NOR2_X1 XNOR_1_3_NUM30 (.ZN (XNOR_1_3_NUM30_OUT), .A1 (XNOR_1_1_NUM30_OUT), .A2 (XNOR_1_2_NUM30_OUT));
      NOR2_X1 XNOR_1_4_NUM30 (.ZN (XNOR_1_4_NUM30_OUT), .A1 (N41), .A2 (N57));
      NOR2_X1 XNOR_1_5_NUM30 (.ZN (N279), .A1 (XNOR_1_3_NUM30_OUT), .A2 (XNOR_1_4_NUM30_OUT));
      wire XNOR_1_1_NUM31_OUT, XNOR_1_2_NUM31_OUT, XNOR_1_3_NUM31_OUT, XNOR_1_4_NUM31_OUT;
      NOR2_X1 XNOR_1_1_NUM31 (.ZN (XNOR_1_1_NUM31_OUT), .A1 (N13), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM31 (.ZN (XNOR_1_2_NUM31_OUT), .A1 (GND), .A2 (N29));
      NOR2_X1 XNOR_1_3_NUM31 (.ZN (XNOR_1_3_NUM31_OUT), .A1 (XNOR_1_1_NUM31_OUT), .A2 (XNOR_1_2_NUM31_OUT));
      NOR2_X1 XNOR_1_4_NUM31 (.ZN (XNOR_1_4_NUM31_OUT), .A1 (N13), .A2 (N29));
      NOR2_X1 XNOR_1_5_NUM31 (.ZN (N280), .A1 (XNOR_1_3_NUM31_OUT), .A2 (XNOR_1_4_NUM31_OUT));
      wire XNOR_1_1_NUM32_OUT, XNOR_1_2_NUM32_OUT, XNOR_1_3_NUM32_OUT, XNOR_1_4_NUM32_OUT;
      NOR2_X1 XNOR_1_1_NUM32 (.ZN (XNOR_1_1_NUM32_OUT), .A1 (N45), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM32 (.ZN (XNOR_1_2_NUM32_OUT), .A1 (GND), .A2 (N61));
      NOR2_X1 XNOR_1_3_NUM32 (.ZN (XNOR_1_3_NUM32_OUT), .A1 (XNOR_1_1_NUM32_OUT), .A2 (XNOR_1_2_NUM32_OUT));
      NOR2_X1 XNOR_1_4_NUM32 (.ZN (XNOR_1_4_NUM32_OUT), .A1 (N45), .A2 (N61));
      NOR2_X1 XNOR_1_5_NUM32 (.ZN (N281), .A1 (XNOR_1_3_NUM32_OUT), .A2 (XNOR_1_4_NUM32_OUT));
      wire XNOR_1_1_NUM33_OUT, XNOR_1_2_NUM33_OUT, XNOR_1_3_NUM33_OUT, XNOR_1_4_NUM33_OUT;
      NOR2_X1 XNOR_1_1_NUM33 (.ZN (XNOR_1_1_NUM33_OUT), .A1 (N65), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM33 (.ZN (XNOR_1_2_NUM33_OUT), .A1 (GND), .A2 (N81));
      NOR2_X1 XNOR_1_3_NUM33 (.ZN (XNOR_1_3_NUM33_OUT), .A1 (XNOR_1_1_NUM33_OUT), .A2 (XNOR_1_2_NUM33_OUT));
      NOR2_X1 XNOR_1_4_NUM33 (.ZN (XNOR_1_4_NUM33_OUT), .A1 (N65), .A2 (N81));
      NOR2_X1 XNOR_1_5_NUM33 (.ZN (N282), .A1 (XNOR_1_3_NUM33_OUT), .A2 (XNOR_1_4_NUM33_OUT));
      wire XNOR_1_1_NUM34_OUT, XNOR_1_2_NUM34_OUT, XNOR_1_3_NUM34_OUT, XNOR_1_4_NUM34_OUT;
      NOR2_X1 XNOR_1_1_NUM34 (.ZN (XNOR_1_1_NUM34_OUT), .A1 (N97), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM34 (.ZN (XNOR_1_2_NUM34_OUT), .A1 (GND), .A2 (N113));
      NOR2_X1 XNOR_1_3_NUM34 (.ZN (XNOR_1_3_NUM34_OUT), .A1 (XNOR_1_1_NUM34_OUT), .A2 (XNOR_1_2_NUM34_OUT));
      NOR2_X1 XNOR_1_4_NUM34 (.ZN (XNOR_1_4_NUM34_OUT), .A1 (N97), .A2 (N113));
      NOR2_X1 XNOR_1_5_NUM34 (.ZN (N283), .A1 (XNOR_1_3_NUM34_OUT), .A2 (XNOR_1_4_NUM34_OUT));
      wire XNOR_1_1_NUM35_OUT, XNOR_1_2_NUM35_OUT, XNOR_1_3_NUM35_OUT, XNOR_1_4_NUM35_OUT;
      NOR2_X1 XNOR_1_1_NUM35 (.ZN (XNOR_1_1_NUM35_OUT), .A1 (N69), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM35 (.ZN (XNOR_1_2_NUM35_OUT), .A1 (GND), .A2 (N85));
      NOR2_X1 XNOR_1_3_NUM35 (.ZN (XNOR_1_3_NUM35_OUT), .A1 (XNOR_1_1_NUM35_OUT), .A2 (XNOR_1_2_NUM35_OUT));
      NOR2_X1 XNOR_1_4_NUM35 (.ZN (XNOR_1_4_NUM35_OUT), .A1 (N69), .A2 (N85));
      NOR2_X1 XNOR_1_5_NUM35 (.ZN (N284), .A1 (XNOR_1_3_NUM35_OUT), .A2 (XNOR_1_4_NUM35_OUT));
      wire XNOR_1_1_NUM36_OUT, XNOR_1_2_NUM36_OUT, XNOR_1_3_NUM36_OUT, XNOR_1_4_NUM36_OUT;
      NOR2_X1 XNOR_1_1_NUM36 (.ZN (XNOR_1_1_NUM36_OUT), .A1 (N101), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM36 (.ZN (XNOR_1_2_NUM36_OUT), .A1 (GND), .A2 (N117));
      NOR2_X1 XNOR_1_3_NUM36 (.ZN (XNOR_1_3_NUM36_OUT), .A1 (XNOR_1_1_NUM36_OUT), .A2 (XNOR_1_2_NUM36_OUT));
      NOR2_X1 XNOR_1_4_NUM36 (.ZN (XNOR_1_4_NUM36_OUT), .A1 (N101), .A2 (N117));
      NOR2_X1 XNOR_1_5_NUM36 (.ZN (N285), .A1 (XNOR_1_3_NUM36_OUT), .A2 (XNOR_1_4_NUM36_OUT));
      wire XNOR_1_1_NUM37_OUT, XNOR_1_2_NUM37_OUT, XNOR_1_3_NUM37_OUT, XNOR_1_4_NUM37_OUT;
      NOR2_X1 XNOR_1_1_NUM37 (.ZN (XNOR_1_1_NUM37_OUT), .A1 (N73), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM37 (.ZN (XNOR_1_2_NUM37_OUT), .A1 (GND), .A2 (N89));
      NOR2_X1 XNOR_1_3_NUM37 (.ZN (XNOR_1_3_NUM37_OUT), .A1 (XNOR_1_1_NUM37_OUT), .A2 (XNOR_1_2_NUM37_OUT));
      NOR2_X1 XNOR_1_4_NUM37 (.ZN (XNOR_1_4_NUM37_OUT), .A1 (N73), .A2 (N89));
      NOR2_X1 XNOR_1_5_NUM37 (.ZN (N286), .A1 (XNOR_1_3_NUM37_OUT), .A2 (XNOR_1_4_NUM37_OUT));
      wire XNOR_1_1_NUM38_OUT, XNOR_1_2_NUM38_OUT, XNOR_1_3_NUM38_OUT, XNOR_1_4_NUM38_OUT;
      NOR2_X1 XNOR_1_1_NUM38 (.ZN (XNOR_1_1_NUM38_OUT), .A1 (N105), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM38 (.ZN (XNOR_1_2_NUM38_OUT), .A1 (GND), .A2 (N121));
      NOR2_X1 XNOR_1_3_NUM38 (.ZN (XNOR_1_3_NUM38_OUT), .A1 (XNOR_1_1_NUM38_OUT), .A2 (XNOR_1_2_NUM38_OUT));
      NOR2_X1 XNOR_1_4_NUM38 (.ZN (XNOR_1_4_NUM38_OUT), .A1 (N105), .A2 (N121));
      NOR2_X1 XNOR_1_5_NUM38 (.ZN (N287), .A1 (XNOR_1_3_NUM38_OUT), .A2 (XNOR_1_4_NUM38_OUT));
      wire XNOR_1_1_NUM39_OUT, XNOR_1_2_NUM39_OUT, XNOR_1_3_NUM39_OUT, XNOR_1_4_NUM39_OUT;
      NOR2_X1 XNOR_1_1_NUM39 (.ZN (XNOR_1_1_NUM39_OUT), .A1 (N77), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM39 (.ZN (XNOR_1_2_NUM39_OUT), .A1 (GND), .A2 (N93));
      NOR2_X1 XNOR_1_3_NUM39 (.ZN (XNOR_1_3_NUM39_OUT), .A1 (XNOR_1_1_NUM39_OUT), .A2 (XNOR_1_2_NUM39_OUT));
      NOR2_X1 XNOR_1_4_NUM39 (.ZN (XNOR_1_4_NUM39_OUT), .A1 (N77), .A2 (N93));
      NOR2_X1 XNOR_1_5_NUM39 (.ZN (N288), .A1 (XNOR_1_3_NUM39_OUT), .A2 (XNOR_1_4_NUM39_OUT));
      wire XNOR_1_1_NUM40_OUT, XNOR_1_2_NUM40_OUT, XNOR_1_3_NUM40_OUT, XNOR_1_4_NUM40_OUT;
      NOR2_X1 XNOR_1_1_NUM40 (.ZN (XNOR_1_1_NUM40_OUT), .A1 (N109), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM40 (.ZN (XNOR_1_2_NUM40_OUT), .A1 (GND), .A2 (N125));
      NOR2_X1 XNOR_1_3_NUM40 (.ZN (XNOR_1_3_NUM40_OUT), .A1 (XNOR_1_1_NUM40_OUT), .A2 (XNOR_1_2_NUM40_OUT));
      NOR2_X1 XNOR_1_4_NUM40 (.ZN (XNOR_1_4_NUM40_OUT), .A1 (N109), .A2 (N125));
      NOR2_X1 XNOR_1_5_NUM40 (.ZN (N289), .A1 (XNOR_1_3_NUM40_OUT), .A2 (XNOR_1_4_NUM40_OUT));
      wire XNOR_1_1_NUM41_OUT, XNOR_1_2_NUM41_OUT, XNOR_1_3_NUM41_OUT, XNOR_1_4_NUM41_OUT;
      NOR2_X1 XNOR_1_1_NUM41 (.ZN (XNOR_1_1_NUM41_OUT), .A1 (N250), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM41 (.ZN (XNOR_1_2_NUM41_OUT), .A1 (GND), .A2 (N251));
      NOR2_X1 XNOR_1_3_NUM41 (.ZN (XNOR_1_3_NUM41_OUT), .A1 (XNOR_1_1_NUM41_OUT), .A2 (XNOR_1_2_NUM41_OUT));
      NOR2_X1 XNOR_1_4_NUM41 (.ZN (XNOR_1_4_NUM41_OUT), .A1 (N250), .A2 (N251));
      NOR2_X1 XNOR_1_5_NUM41 (.ZN (N290), .A1 (XNOR_1_3_NUM41_OUT), .A2 (XNOR_1_4_NUM41_OUT));
      wire XNOR_1_1_NUM42_OUT, XNOR_1_2_NUM42_OUT, XNOR_1_3_NUM42_OUT, XNOR_1_4_NUM42_OUT;
      NOR2_X1 XNOR_1_1_NUM42 (.ZN (XNOR_1_1_NUM42_OUT), .A1 (N252), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM42 (.ZN (XNOR_1_2_NUM42_OUT), .A1 (GND), .A2 (N253));
      NOR2_X1 XNOR_1_3_NUM42 (.ZN (XNOR_1_3_NUM42_OUT), .A1 (XNOR_1_1_NUM42_OUT), .A2 (XNOR_1_2_NUM42_OUT));
      NOR2_X1 XNOR_1_4_NUM42 (.ZN (XNOR_1_4_NUM42_OUT), .A1 (N252), .A2 (N253));
      NOR2_X1 XNOR_1_5_NUM42 (.ZN (N293), .A1 (XNOR_1_3_NUM42_OUT), .A2 (XNOR_1_4_NUM42_OUT));
      wire XNOR_1_1_NUM43_OUT, XNOR_1_2_NUM43_OUT, XNOR_1_3_NUM43_OUT, XNOR_1_4_NUM43_OUT;
      NOR2_X1 XNOR_1_1_NUM43 (.ZN (XNOR_1_1_NUM43_OUT), .A1 (N254), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM43 (.ZN (XNOR_1_2_NUM43_OUT), .A1 (GND), .A2 (N255));
      NOR2_X1 XNOR_1_3_NUM43 (.ZN (XNOR_1_3_NUM43_OUT), .A1 (XNOR_1_1_NUM43_OUT), .A2 (XNOR_1_2_NUM43_OUT));
      NOR2_X1 XNOR_1_4_NUM43 (.ZN (XNOR_1_4_NUM43_OUT), .A1 (N254), .A2 (N255));
      NOR2_X1 XNOR_1_5_NUM43 (.ZN (N296), .A1 (XNOR_1_3_NUM43_OUT), .A2 (XNOR_1_4_NUM43_OUT));
      wire XNOR_1_1_NUM44_OUT, XNOR_1_2_NUM44_OUT, XNOR_1_3_NUM44_OUT, XNOR_1_4_NUM44_OUT;
      NOR2_X1 XNOR_1_1_NUM44 (.ZN (XNOR_1_1_NUM44_OUT), .A1 (N256), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM44 (.ZN (XNOR_1_2_NUM44_OUT), .A1 (GND), .A2 (N257));
      NOR2_X1 XNOR_1_3_NUM44 (.ZN (XNOR_1_3_NUM44_OUT), .A1 (XNOR_1_1_NUM44_OUT), .A2 (XNOR_1_2_NUM44_OUT));
      NOR2_X1 XNOR_1_4_NUM44 (.ZN (XNOR_1_4_NUM44_OUT), .A1 (N256), .A2 (N257));
      NOR2_X1 XNOR_1_5_NUM44 (.ZN (N299), .A1 (XNOR_1_3_NUM44_OUT), .A2 (XNOR_1_4_NUM44_OUT));
      wire XNOR_1_1_NUM45_OUT, XNOR_1_2_NUM45_OUT, XNOR_1_3_NUM45_OUT, XNOR_1_4_NUM45_OUT;
      NOR2_X1 XNOR_1_1_NUM45 (.ZN (XNOR_1_1_NUM45_OUT), .A1 (N258), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM45 (.ZN (XNOR_1_2_NUM45_OUT), .A1 (GND), .A2 (N259));
      NOR2_X1 XNOR_1_3_NUM45 (.ZN (XNOR_1_3_NUM45_OUT), .A1 (XNOR_1_1_NUM45_OUT), .A2 (XNOR_1_2_NUM45_OUT));
      NOR2_X1 XNOR_1_4_NUM45 (.ZN (XNOR_1_4_NUM45_OUT), .A1 (N258), .A2 (N259));
      NOR2_X1 XNOR_1_5_NUM45 (.ZN (N302), .A1 (XNOR_1_3_NUM45_OUT), .A2 (XNOR_1_4_NUM45_OUT));
      wire XNOR_1_1_NUM46_OUT, XNOR_1_2_NUM46_OUT, XNOR_1_3_NUM46_OUT, XNOR_1_4_NUM46_OUT;
      NOR2_X1 XNOR_1_1_NUM46 (.ZN (XNOR_1_1_NUM46_OUT), .A1 (N260), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM46 (.ZN (XNOR_1_2_NUM46_OUT), .A1 (GND), .A2 (N261));
      NOR2_X1 XNOR_1_3_NUM46 (.ZN (XNOR_1_3_NUM46_OUT), .A1 (XNOR_1_1_NUM46_OUT), .A2 (XNOR_1_2_NUM46_OUT));
      NOR2_X1 XNOR_1_4_NUM46 (.ZN (XNOR_1_4_NUM46_OUT), .A1 (N260), .A2 (N261));
      NOR2_X1 XNOR_1_5_NUM46 (.ZN (N305), .A1 (XNOR_1_3_NUM46_OUT), .A2 (XNOR_1_4_NUM46_OUT));
      wire XNOR_1_1_NUM47_OUT, XNOR_1_2_NUM47_OUT, XNOR_1_3_NUM47_OUT, XNOR_1_4_NUM47_OUT;
      NOR2_X1 XNOR_1_1_NUM47 (.ZN (XNOR_1_1_NUM47_OUT), .A1 (N262), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM47 (.ZN (XNOR_1_2_NUM47_OUT), .A1 (GND), .A2 (N263));
      NOR2_X1 XNOR_1_3_NUM47 (.ZN (XNOR_1_3_NUM47_OUT), .A1 (XNOR_1_1_NUM47_OUT), .A2 (XNOR_1_2_NUM47_OUT));
      NOR2_X1 XNOR_1_4_NUM47 (.ZN (XNOR_1_4_NUM47_OUT), .A1 (N262), .A2 (N263));
      NOR2_X1 XNOR_1_5_NUM47 (.ZN (N308), .A1 (XNOR_1_3_NUM47_OUT), .A2 (XNOR_1_4_NUM47_OUT));
      wire XNOR_1_1_NUM48_OUT, XNOR_1_2_NUM48_OUT, XNOR_1_3_NUM48_OUT, XNOR_1_4_NUM48_OUT;
      NOR2_X1 XNOR_1_1_NUM48 (.ZN (XNOR_1_1_NUM48_OUT), .A1 (N264), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM48 (.ZN (XNOR_1_2_NUM48_OUT), .A1 (GND), .A2 (N265));
      NOR2_X1 XNOR_1_3_NUM48 (.ZN (XNOR_1_3_NUM48_OUT), .A1 (XNOR_1_1_NUM48_OUT), .A2 (XNOR_1_2_NUM48_OUT));
      NOR2_X1 XNOR_1_4_NUM48 (.ZN (XNOR_1_4_NUM48_OUT), .A1 (N264), .A2 (N265));
      NOR2_X1 XNOR_1_5_NUM48 (.ZN (N311), .A1 (XNOR_1_3_NUM48_OUT), .A2 (XNOR_1_4_NUM48_OUT));
      wire XNOR_1_1_NUM49_OUT, XNOR_1_2_NUM49_OUT, XNOR_1_3_NUM49_OUT, XNOR_1_4_NUM49_OUT;
      NOR2_X1 XNOR_1_1_NUM49 (.ZN (XNOR_1_1_NUM49_OUT), .A1 (N274), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM49 (.ZN (XNOR_1_2_NUM49_OUT), .A1 (GND), .A2 (N275));
      NOR2_X1 XNOR_1_3_NUM49 (.ZN (XNOR_1_3_NUM49_OUT), .A1 (XNOR_1_1_NUM49_OUT), .A2 (XNOR_1_2_NUM49_OUT));
      NOR2_X1 XNOR_1_4_NUM49 (.ZN (XNOR_1_4_NUM49_OUT), .A1 (N274), .A2 (N275));
      NOR2_X1 XNOR_1_5_NUM49 (.ZN (N314), .A1 (XNOR_1_3_NUM49_OUT), .A2 (XNOR_1_4_NUM49_OUT));
      wire XNOR_1_1_NUM50_OUT, XNOR_1_2_NUM50_OUT, XNOR_1_3_NUM50_OUT, XNOR_1_4_NUM50_OUT;
      NOR2_X1 XNOR_1_1_NUM50 (.ZN (XNOR_1_1_NUM50_OUT), .A1 (N276), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM50 (.ZN (XNOR_1_2_NUM50_OUT), .A1 (GND), .A2 (N277));
      NOR2_X1 XNOR_1_3_NUM50 (.ZN (XNOR_1_3_NUM50_OUT), .A1 (XNOR_1_1_NUM50_OUT), .A2 (XNOR_1_2_NUM50_OUT));
      NOR2_X1 XNOR_1_4_NUM50 (.ZN (XNOR_1_4_NUM50_OUT), .A1 (N276), .A2 (N277));
      NOR2_X1 XNOR_1_5_NUM50 (.ZN (N315), .A1 (XNOR_1_3_NUM50_OUT), .A2 (XNOR_1_4_NUM50_OUT));
      wire XNOR_1_1_NUM51_OUT, XNOR_1_2_NUM51_OUT, XNOR_1_3_NUM51_OUT, XNOR_1_4_NUM51_OUT;
      NOR2_X1 XNOR_1_1_NUM51 (.ZN (XNOR_1_1_NUM51_OUT), .A1 (N278), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM51 (.ZN (XNOR_1_2_NUM51_OUT), .A1 (GND), .A2 (N279));
      NOR2_X1 XNOR_1_3_NUM51 (.ZN (XNOR_1_3_NUM51_OUT), .A1 (XNOR_1_1_NUM51_OUT), .A2 (XNOR_1_2_NUM51_OUT));
      NOR2_X1 XNOR_1_4_NUM51 (.ZN (XNOR_1_4_NUM51_OUT), .A1 (N278), .A2 (N279));
      NOR2_X1 XNOR_1_5_NUM51 (.ZN (N316), .A1 (XNOR_1_3_NUM51_OUT), .A2 (XNOR_1_4_NUM51_OUT));
      wire XNOR_1_1_NUM52_OUT, XNOR_1_2_NUM52_OUT, XNOR_1_3_NUM52_OUT, XNOR_1_4_NUM52_OUT;
      NOR2_X1 XNOR_1_1_NUM52 (.ZN (XNOR_1_1_NUM52_OUT), .A1 (N280), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM52 (.ZN (XNOR_1_2_NUM52_OUT), .A1 (GND), .A2 (N281));
      NOR2_X1 XNOR_1_3_NUM52 (.ZN (XNOR_1_3_NUM52_OUT), .A1 (XNOR_1_1_NUM52_OUT), .A2 (XNOR_1_2_NUM52_OUT));
      NOR2_X1 XNOR_1_4_NUM52 (.ZN (XNOR_1_4_NUM52_OUT), .A1 (N280), .A2 (N281));
      NOR2_X1 XNOR_1_5_NUM52 (.ZN (N317), .A1 (XNOR_1_3_NUM52_OUT), .A2 (XNOR_1_4_NUM52_OUT));
      wire XNOR_1_1_NUM53_OUT, XNOR_1_2_NUM53_OUT, XNOR_1_3_NUM53_OUT, XNOR_1_4_NUM53_OUT;
      NOR2_X1 XNOR_1_1_NUM53 (.ZN (XNOR_1_1_NUM53_OUT), .A1 (N282), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM53 (.ZN (XNOR_1_2_NUM53_OUT), .A1 (GND), .A2 (N283));
      NOR2_X1 XNOR_1_3_NUM53 (.ZN (XNOR_1_3_NUM53_OUT), .A1 (XNOR_1_1_NUM53_OUT), .A2 (XNOR_1_2_NUM53_OUT));
      NOR2_X1 XNOR_1_4_NUM53 (.ZN (XNOR_1_4_NUM53_OUT), .A1 (N282), .A2 (N283));
      NOR2_X1 XNOR_1_5_NUM53 (.ZN (N318), .A1 (XNOR_1_3_NUM53_OUT), .A2 (XNOR_1_4_NUM53_OUT));
      wire XNOR_1_1_NUM54_OUT, XNOR_1_2_NUM54_OUT, XNOR_1_3_NUM54_OUT, XNOR_1_4_NUM54_OUT;
      NOR2_X1 XNOR_1_1_NUM54 (.ZN (XNOR_1_1_NUM54_OUT), .A1 (N284), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM54 (.ZN (XNOR_1_2_NUM54_OUT), .A1 (GND), .A2 (N285));
      NOR2_X1 XNOR_1_3_NUM54 (.ZN (XNOR_1_3_NUM54_OUT), .A1 (XNOR_1_1_NUM54_OUT), .A2 (XNOR_1_2_NUM54_OUT));
      NOR2_X1 XNOR_1_4_NUM54 (.ZN (XNOR_1_4_NUM54_OUT), .A1 (N284), .A2 (N285));
      NOR2_X1 XNOR_1_5_NUM54 (.ZN (N319), .A1 (XNOR_1_3_NUM54_OUT), .A2 (XNOR_1_4_NUM54_OUT));
      wire XNOR_1_1_NUM55_OUT, XNOR_1_2_NUM55_OUT, XNOR_1_3_NUM55_OUT, XNOR_1_4_NUM55_OUT;
      NOR2_X1 XNOR_1_1_NUM55 (.ZN (XNOR_1_1_NUM55_OUT), .A1 (N286), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM55 (.ZN (XNOR_1_2_NUM55_OUT), .A1 (GND), .A2 (N287));
      NOR2_X1 XNOR_1_3_NUM55 (.ZN (XNOR_1_3_NUM55_OUT), .A1 (XNOR_1_1_NUM55_OUT), .A2 (XNOR_1_2_NUM55_OUT));
      NOR2_X1 XNOR_1_4_NUM55 (.ZN (XNOR_1_4_NUM55_OUT), .A1 (N286), .A2 (N287));
      NOR2_X1 XNOR_1_5_NUM55 (.ZN (N320), .A1 (XNOR_1_3_NUM55_OUT), .A2 (XNOR_1_4_NUM55_OUT));
      wire XNOR_1_1_NUM56_OUT, XNOR_1_2_NUM56_OUT, XNOR_1_3_NUM56_OUT, XNOR_1_4_NUM56_OUT;
      NOR2_X1 XNOR_1_1_NUM56 (.ZN (XNOR_1_1_NUM56_OUT), .A1 (N288), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM56 (.ZN (XNOR_1_2_NUM56_OUT), .A1 (GND), .A2 (N289));
      NOR2_X1 XNOR_1_3_NUM56 (.ZN (XNOR_1_3_NUM56_OUT), .A1 (XNOR_1_1_NUM56_OUT), .A2 (XNOR_1_2_NUM56_OUT));
      NOR2_X1 XNOR_1_4_NUM56 (.ZN (XNOR_1_4_NUM56_OUT), .A1 (N288), .A2 (N289));
      NOR2_X1 XNOR_1_5_NUM56 (.ZN (N321), .A1 (XNOR_1_3_NUM56_OUT), .A2 (XNOR_1_4_NUM56_OUT));
      wire XNOR_1_1_NUM57_OUT, XNOR_1_2_NUM57_OUT, XNOR_1_3_NUM57_OUT, XNOR_1_4_NUM57_OUT;
      NOR2_X1 XNOR_1_1_NUM57 (.ZN (XNOR_1_1_NUM57_OUT), .A1 (N290), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM57 (.ZN (XNOR_1_2_NUM57_OUT), .A1 (GND), .A2 (N293));
      NOR2_X1 XNOR_1_3_NUM57 (.ZN (XNOR_1_3_NUM57_OUT), .A1 (XNOR_1_1_NUM57_OUT), .A2 (XNOR_1_2_NUM57_OUT));
      NOR2_X1 XNOR_1_4_NUM57 (.ZN (XNOR_1_4_NUM57_OUT), .A1 (N290), .A2 (N293));
      NOR2_X1 XNOR_1_5_NUM57 (.ZN (N338), .A1 (XNOR_1_3_NUM57_OUT), .A2 (XNOR_1_4_NUM57_OUT));
      wire XNOR_1_1_NUM58_OUT, XNOR_1_2_NUM58_OUT, XNOR_1_3_NUM58_OUT, XNOR_1_4_NUM58_OUT;
      NOR2_X1 XNOR_1_1_NUM58 (.ZN (XNOR_1_1_NUM58_OUT), .A1 (N296), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM58 (.ZN (XNOR_1_2_NUM58_OUT), .A1 (GND), .A2 (N299));
      NOR2_X1 XNOR_1_3_NUM58 (.ZN (XNOR_1_3_NUM58_OUT), .A1 (XNOR_1_1_NUM58_OUT), .A2 (XNOR_1_2_NUM58_OUT));
      NOR2_X1 XNOR_1_4_NUM58 (.ZN (XNOR_1_4_NUM58_OUT), .A1 (N296), .A2 (N299));
      NOR2_X1 XNOR_1_5_NUM58 (.ZN (N339), .A1 (XNOR_1_3_NUM58_OUT), .A2 (XNOR_1_4_NUM58_OUT));
      wire XNOR_1_1_NUM59_OUT, XNOR_1_2_NUM59_OUT, XNOR_1_3_NUM59_OUT, XNOR_1_4_NUM59_OUT;
      NOR2_X1 XNOR_1_1_NUM59 (.ZN (XNOR_1_1_NUM59_OUT), .A1 (N290), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM59 (.ZN (XNOR_1_2_NUM59_OUT), .A1 (GND), .A2 (N296));
      NOR2_X1 XNOR_1_3_NUM59 (.ZN (XNOR_1_3_NUM59_OUT), .A1 (XNOR_1_1_NUM59_OUT), .A2 (XNOR_1_2_NUM59_OUT));
      NOR2_X1 XNOR_1_4_NUM59 (.ZN (XNOR_1_4_NUM59_OUT), .A1 (N290), .A2 (N296));
      NOR2_X1 XNOR_1_5_NUM59 (.ZN (N340), .A1 (XNOR_1_3_NUM59_OUT), .A2 (XNOR_1_4_NUM59_OUT));
      wire XNOR_1_1_NUM60_OUT, XNOR_1_2_NUM60_OUT, XNOR_1_3_NUM60_OUT, XNOR_1_4_NUM60_OUT;
      NOR2_X1 XNOR_1_1_NUM60 (.ZN (XNOR_1_1_NUM60_OUT), .A1 (N293), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM60 (.ZN (XNOR_1_2_NUM60_OUT), .A1 (GND), .A2 (N299));
      NOR2_X1 XNOR_1_3_NUM60 (.ZN (XNOR_1_3_NUM60_OUT), .A1 (XNOR_1_1_NUM60_OUT), .A2 (XNOR_1_2_NUM60_OUT));
      NOR2_X1 XNOR_1_4_NUM60 (.ZN (XNOR_1_4_NUM60_OUT), .A1 (N293), .A2 (N299));
      NOR2_X1 XNOR_1_5_NUM60 (.ZN (N341), .A1 (XNOR_1_3_NUM60_OUT), .A2 (XNOR_1_4_NUM60_OUT));
      wire XNOR_1_1_NUM61_OUT, XNOR_1_2_NUM61_OUT, XNOR_1_3_NUM61_OUT, XNOR_1_4_NUM61_OUT;
      NOR2_X1 XNOR_1_1_NUM61 (.ZN (XNOR_1_1_NUM61_OUT), .A1 (N302), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM61 (.ZN (XNOR_1_2_NUM61_OUT), .A1 (GND), .A2 (N305));
      NOR2_X1 XNOR_1_3_NUM61 (.ZN (XNOR_1_3_NUM61_OUT), .A1 (XNOR_1_1_NUM61_OUT), .A2 (XNOR_1_2_NUM61_OUT));
      NOR2_X1 XNOR_1_4_NUM61 (.ZN (XNOR_1_4_NUM61_OUT), .A1 (N302), .A2 (N305));
      NOR2_X1 XNOR_1_5_NUM61 (.ZN (N342), .A1 (XNOR_1_3_NUM61_OUT), .A2 (XNOR_1_4_NUM61_OUT));
      wire XNOR_1_1_NUM62_OUT, XNOR_1_2_NUM62_OUT, XNOR_1_3_NUM62_OUT, XNOR_1_4_NUM62_OUT;
      NOR2_X1 XNOR_1_1_NUM62 (.ZN (XNOR_1_1_NUM62_OUT), .A1 (N308), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM62 (.ZN (XNOR_1_2_NUM62_OUT), .A1 (GND), .A2 (N311));
      NOR2_X1 XNOR_1_3_NUM62 (.ZN (XNOR_1_3_NUM62_OUT), .A1 (XNOR_1_1_NUM62_OUT), .A2 (XNOR_1_2_NUM62_OUT));
      NOR2_X1 XNOR_1_4_NUM62 (.ZN (XNOR_1_4_NUM62_OUT), .A1 (N308), .A2 (N311));
      NOR2_X1 XNOR_1_5_NUM62 (.ZN (N343), .A1 (XNOR_1_3_NUM62_OUT), .A2 (XNOR_1_4_NUM62_OUT));
      wire XNOR_1_1_NUM63_OUT, XNOR_1_2_NUM63_OUT, XNOR_1_3_NUM63_OUT, XNOR_1_4_NUM63_OUT;
      NOR2_X1 XNOR_1_1_NUM63 (.ZN (XNOR_1_1_NUM63_OUT), .A1 (N302), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM63 (.ZN (XNOR_1_2_NUM63_OUT), .A1 (GND), .A2 (N308));
      NOR2_X1 XNOR_1_3_NUM63 (.ZN (XNOR_1_3_NUM63_OUT), .A1 (XNOR_1_1_NUM63_OUT), .A2 (XNOR_1_2_NUM63_OUT));
      NOR2_X1 XNOR_1_4_NUM63 (.ZN (XNOR_1_4_NUM63_OUT), .A1 (N302), .A2 (N308));
      NOR2_X1 XNOR_1_5_NUM63 (.ZN (N344), .A1 (XNOR_1_3_NUM63_OUT), .A2 (XNOR_1_4_NUM63_OUT));
      wire XNOR_1_1_NUM64_OUT, XNOR_1_2_NUM64_OUT, XNOR_1_3_NUM64_OUT, XNOR_1_4_NUM64_OUT;
      NOR2_X1 XNOR_1_1_NUM64 (.ZN (XNOR_1_1_NUM64_OUT), .A1 (N305), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM64 (.ZN (XNOR_1_2_NUM64_OUT), .A1 (GND), .A2 (N311));
      NOR2_X1 XNOR_1_3_NUM64 (.ZN (XNOR_1_3_NUM64_OUT), .A1 (XNOR_1_1_NUM64_OUT), .A2 (XNOR_1_2_NUM64_OUT));
      NOR2_X1 XNOR_1_4_NUM64 (.ZN (XNOR_1_4_NUM64_OUT), .A1 (N305), .A2 (N311));
      NOR2_X1 XNOR_1_5_NUM64 (.ZN (N345), .A1 (XNOR_1_3_NUM64_OUT), .A2 (XNOR_1_4_NUM64_OUT));
      wire XNOR_1_1_NUM65_OUT, XNOR_1_2_NUM65_OUT, XNOR_1_3_NUM65_OUT, XNOR_1_4_NUM65_OUT;
      NOR2_X1 XNOR_1_1_NUM65 (.ZN (XNOR_1_1_NUM65_OUT), .A1 (N266), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM65 (.ZN (XNOR_1_2_NUM65_OUT), .A1 (GND), .A2 (N342));
      NOR2_X1 XNOR_1_3_NUM65 (.ZN (XNOR_1_3_NUM65_OUT), .A1 (XNOR_1_1_NUM65_OUT), .A2 (XNOR_1_2_NUM65_OUT));
      NOR2_X1 XNOR_1_4_NUM65 (.ZN (XNOR_1_4_NUM65_OUT), .A1 (N266), .A2 (N342));
      NOR2_X1 XNOR_1_5_NUM65 (.ZN (N346), .A1 (XNOR_1_3_NUM65_OUT), .A2 (XNOR_1_4_NUM65_OUT));
      wire XNOR_1_1_NUM66_OUT, XNOR_1_2_NUM66_OUT, XNOR_1_3_NUM66_OUT, XNOR_1_4_NUM66_OUT;
      NOR2_X1 XNOR_1_1_NUM66 (.ZN (XNOR_1_1_NUM66_OUT), .A1 (N267), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM66 (.ZN (XNOR_1_2_NUM66_OUT), .A1 (GND), .A2 (N343));
      NOR2_X1 XNOR_1_3_NUM66 (.ZN (XNOR_1_3_NUM66_OUT), .A1 (XNOR_1_1_NUM66_OUT), .A2 (XNOR_1_2_NUM66_OUT));
      NOR2_X1 XNOR_1_4_NUM66 (.ZN (XNOR_1_4_NUM66_OUT), .A1 (N267), .A2 (N343));
      NOR2_X1 XNOR_1_5_NUM66 (.ZN (N347), .A1 (XNOR_1_3_NUM66_OUT), .A2 (XNOR_1_4_NUM66_OUT));
      wire XNOR_1_1_NUM67_OUT, XNOR_1_2_NUM67_OUT, XNOR_1_3_NUM67_OUT, XNOR_1_4_NUM67_OUT;
      NOR2_X1 XNOR_1_1_NUM67 (.ZN (XNOR_1_1_NUM67_OUT), .A1 (N268), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM67 (.ZN (XNOR_1_2_NUM67_OUT), .A1 (GND), .A2 (N344));
      NOR2_X1 XNOR_1_3_NUM67 (.ZN (XNOR_1_3_NUM67_OUT), .A1 (XNOR_1_1_NUM67_OUT), .A2 (XNOR_1_2_NUM67_OUT));
      NOR2_X1 XNOR_1_4_NUM67 (.ZN (XNOR_1_4_NUM67_OUT), .A1 (N268), .A2 (N344));
      NOR2_X1 XNOR_1_5_NUM67 (.ZN (N348), .A1 (XNOR_1_3_NUM67_OUT), .A2 (XNOR_1_4_NUM67_OUT));
      wire XNOR_1_1_NUM68_OUT, XNOR_1_2_NUM68_OUT, XNOR_1_3_NUM68_OUT, XNOR_1_4_NUM68_OUT;
      NOR2_X1 XNOR_1_1_NUM68 (.ZN (XNOR_1_1_NUM68_OUT), .A1 (N269), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM68 (.ZN (XNOR_1_2_NUM68_OUT), .A1 (GND), .A2 (N345));
      NOR2_X1 XNOR_1_3_NUM68 (.ZN (XNOR_1_3_NUM68_OUT), .A1 (XNOR_1_1_NUM68_OUT), .A2 (XNOR_1_2_NUM68_OUT));
      NOR2_X1 XNOR_1_4_NUM68 (.ZN (XNOR_1_4_NUM68_OUT), .A1 (N269), .A2 (N345));
      NOR2_X1 XNOR_1_5_NUM68 (.ZN (N349), .A1 (XNOR_1_3_NUM68_OUT), .A2 (XNOR_1_4_NUM68_OUT));
      wire XNOR_1_1_NUM69_OUT, XNOR_1_2_NUM69_OUT, XNOR_1_3_NUM69_OUT, XNOR_1_4_NUM69_OUT;
      NOR2_X1 XNOR_1_1_NUM69 (.ZN (XNOR_1_1_NUM69_OUT), .A1 (N270), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM69 (.ZN (XNOR_1_2_NUM69_OUT), .A1 (GND), .A2 (N338));
      NOR2_X1 XNOR_1_3_NUM69 (.ZN (XNOR_1_3_NUM69_OUT), .A1 (XNOR_1_1_NUM69_OUT), .A2 (XNOR_1_2_NUM69_OUT));
      NOR2_X1 XNOR_1_4_NUM69 (.ZN (XNOR_1_4_NUM69_OUT), .A1 (N270), .A2 (N338));
      NOR2_X1 XNOR_1_5_NUM69 (.ZN (N350), .A1 (XNOR_1_3_NUM69_OUT), .A2 (XNOR_1_4_NUM69_OUT));
      wire XNOR_1_1_NUM70_OUT, XNOR_1_2_NUM70_OUT, XNOR_1_3_NUM70_OUT, XNOR_1_4_NUM70_OUT;
      NOR2_X1 XNOR_1_1_NUM70 (.ZN (XNOR_1_1_NUM70_OUT), .A1 (N271), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM70 (.ZN (XNOR_1_2_NUM70_OUT), .A1 (GND), .A2 (N339));
      NOR2_X1 XNOR_1_3_NUM70 (.ZN (XNOR_1_3_NUM70_OUT), .A1 (XNOR_1_1_NUM70_OUT), .A2 (XNOR_1_2_NUM70_OUT));
      NOR2_X1 XNOR_1_4_NUM70 (.ZN (XNOR_1_4_NUM70_OUT), .A1 (N271), .A2 (N339));
      NOR2_X1 XNOR_1_5_NUM70 (.ZN (N351), .A1 (XNOR_1_3_NUM70_OUT), .A2 (XNOR_1_4_NUM70_OUT));
      wire XNOR_1_1_NUM71_OUT, XNOR_1_2_NUM71_OUT, XNOR_1_3_NUM71_OUT, XNOR_1_4_NUM71_OUT;
      NOR2_X1 XNOR_1_1_NUM71 (.ZN (XNOR_1_1_NUM71_OUT), .A1 (N272), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM71 (.ZN (XNOR_1_2_NUM71_OUT), .A1 (GND), .A2 (N340));
      NOR2_X1 XNOR_1_3_NUM71 (.ZN (XNOR_1_3_NUM71_OUT), .A1 (XNOR_1_1_NUM71_OUT), .A2 (XNOR_1_2_NUM71_OUT));
      NOR2_X1 XNOR_1_4_NUM71 (.ZN (XNOR_1_4_NUM71_OUT), .A1 (N272), .A2 (N340));
      NOR2_X1 XNOR_1_5_NUM71 (.ZN (N352), .A1 (XNOR_1_3_NUM71_OUT), .A2 (XNOR_1_4_NUM71_OUT));
      wire XNOR_1_1_NUM72_OUT, XNOR_1_2_NUM72_OUT, XNOR_1_3_NUM72_OUT, XNOR_1_4_NUM72_OUT;
      NOR2_X1 XNOR_1_1_NUM72 (.ZN (XNOR_1_1_NUM72_OUT), .A1 (N273), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM72 (.ZN (XNOR_1_2_NUM72_OUT), .A1 (GND), .A2 (N341));
      NOR2_X1 XNOR_1_3_NUM72 (.ZN (XNOR_1_3_NUM72_OUT), .A1 (XNOR_1_1_NUM72_OUT), .A2 (XNOR_1_2_NUM72_OUT));
      NOR2_X1 XNOR_1_4_NUM72 (.ZN (XNOR_1_4_NUM72_OUT), .A1 (N273), .A2 (N341));
      NOR2_X1 XNOR_1_5_NUM72 (.ZN (N353), .A1 (XNOR_1_3_NUM72_OUT), .A2 (XNOR_1_4_NUM72_OUT));
      wire XNOR_1_1_NUM73_OUT, XNOR_1_2_NUM73_OUT, XNOR_1_3_NUM73_OUT, XNOR_1_4_NUM73_OUT;
      NOR2_X1 XNOR_1_1_NUM73 (.ZN (XNOR_1_1_NUM73_OUT), .A1 (N314), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM73 (.ZN (XNOR_1_2_NUM73_OUT), .A1 (GND), .A2 (N346));
      NOR2_X1 XNOR_1_3_NUM73 (.ZN (XNOR_1_3_NUM73_OUT), .A1 (XNOR_1_1_NUM73_OUT), .A2 (XNOR_1_2_NUM73_OUT));
      NOR2_X1 XNOR_1_4_NUM73 (.ZN (XNOR_1_4_NUM73_OUT), .A1 (N314), .A2 (N346));
      NOR2_X1 XNOR_1_5_NUM73 (.ZN (N354), .A1 (XNOR_1_3_NUM73_OUT), .A2 (XNOR_1_4_NUM73_OUT));
      wire XNOR_1_1_NUM74_OUT, XNOR_1_2_NUM74_OUT, XNOR_1_3_NUM74_OUT, XNOR_1_4_NUM74_OUT;
      NOR2_X1 XNOR_1_1_NUM74 (.ZN (XNOR_1_1_NUM74_OUT), .A1 (N315), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM74 (.ZN (XNOR_1_2_NUM74_OUT), .A1 (GND), .A2 (N347));
      NOR2_X1 XNOR_1_3_NUM74 (.ZN (XNOR_1_3_NUM74_OUT), .A1 (XNOR_1_1_NUM74_OUT), .A2 (XNOR_1_2_NUM74_OUT));
      NOR2_X1 XNOR_1_4_NUM74 (.ZN (XNOR_1_4_NUM74_OUT), .A1 (N315), .A2 (N347));
      NOR2_X1 XNOR_1_5_NUM74 (.ZN (N367), .A1 (XNOR_1_3_NUM74_OUT), .A2 (XNOR_1_4_NUM74_OUT));
      wire XNOR_1_1_NUM75_OUT, XNOR_1_2_NUM75_OUT, XNOR_1_3_NUM75_OUT, XNOR_1_4_NUM75_OUT;
      NOR2_X1 XNOR_1_1_NUM75 (.ZN (XNOR_1_1_NUM75_OUT), .A1 (N316), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM75 (.ZN (XNOR_1_2_NUM75_OUT), .A1 (GND), .A2 (N348));
      NOR2_X1 XNOR_1_3_NUM75 (.ZN (XNOR_1_3_NUM75_OUT), .A1 (XNOR_1_1_NUM75_OUT), .A2 (XNOR_1_2_NUM75_OUT));
      NOR2_X1 XNOR_1_4_NUM75 (.ZN (XNOR_1_4_NUM75_OUT), .A1 (N316), .A2 (N348));
      NOR2_X1 XNOR_1_5_NUM75 (.ZN (N380), .A1 (XNOR_1_3_NUM75_OUT), .A2 (XNOR_1_4_NUM75_OUT));
      wire XNOR_1_1_NUM76_OUT, XNOR_1_2_NUM76_OUT, XNOR_1_3_NUM76_OUT, XNOR_1_4_NUM76_OUT;
      NOR2_X1 XNOR_1_1_NUM76 (.ZN (XNOR_1_1_NUM76_OUT), .A1 (N317), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM76 (.ZN (XNOR_1_2_NUM76_OUT), .A1 (GND), .A2 (N349));
      NOR2_X1 XNOR_1_3_NUM76 (.ZN (XNOR_1_3_NUM76_OUT), .A1 (XNOR_1_1_NUM76_OUT), .A2 (XNOR_1_2_NUM76_OUT));
      NOR2_X1 XNOR_1_4_NUM76 (.ZN (XNOR_1_4_NUM76_OUT), .A1 (N317), .A2 (N349));
      NOR2_X1 XNOR_1_5_NUM76 (.ZN (N393), .A1 (XNOR_1_3_NUM76_OUT), .A2 (XNOR_1_4_NUM76_OUT));
      wire XNOR_1_1_NUM77_OUT, XNOR_1_2_NUM77_OUT, XNOR_1_3_NUM77_OUT, XNOR_1_4_NUM77_OUT;
      NOR2_X1 XNOR_1_1_NUM77 (.ZN (XNOR_1_1_NUM77_OUT), .A1 (N318), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM77 (.ZN (XNOR_1_2_NUM77_OUT), .A1 (GND), .A2 (N350));
      NOR2_X1 XNOR_1_3_NUM77 (.ZN (XNOR_1_3_NUM77_OUT), .A1 (XNOR_1_1_NUM77_OUT), .A2 (XNOR_1_2_NUM77_OUT));
      NOR2_X1 XNOR_1_4_NUM77 (.ZN (XNOR_1_4_NUM77_OUT), .A1 (N318), .A2 (N350));
      NOR2_X1 XNOR_1_5_NUM77 (.ZN (N406), .A1 (XNOR_1_3_NUM77_OUT), .A2 (XNOR_1_4_NUM77_OUT));
      wire XNOR_1_1_NUM78_OUT, XNOR_1_2_NUM78_OUT, XNOR_1_3_NUM78_OUT, XNOR_1_4_NUM78_OUT;
      NOR2_X1 XNOR_1_1_NUM78 (.ZN (XNOR_1_1_NUM78_OUT), .A1 (N319), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM78 (.ZN (XNOR_1_2_NUM78_OUT), .A1 (GND), .A2 (N351));
      NOR2_X1 XNOR_1_3_NUM78 (.ZN (XNOR_1_3_NUM78_OUT), .A1 (XNOR_1_1_NUM78_OUT), .A2 (XNOR_1_2_NUM78_OUT));
      NOR2_X1 XNOR_1_4_NUM78 (.ZN (XNOR_1_4_NUM78_OUT), .A1 (N319), .A2 (N351));
      NOR2_X1 XNOR_1_5_NUM78 (.ZN (N419), .A1 (XNOR_1_3_NUM78_OUT), .A2 (XNOR_1_4_NUM78_OUT));
      wire XNOR_1_1_NUM79_OUT, XNOR_1_2_NUM79_OUT, XNOR_1_3_NUM79_OUT, XNOR_1_4_NUM79_OUT;
      NOR2_X1 XNOR_1_1_NUM79 (.ZN (XNOR_1_1_NUM79_OUT), .A1 (N320), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM79 (.ZN (XNOR_1_2_NUM79_OUT), .A1 (GND), .A2 (N352));
      NOR2_X1 XNOR_1_3_NUM79 (.ZN (XNOR_1_3_NUM79_OUT), .A1 (XNOR_1_1_NUM79_OUT), .A2 (XNOR_1_2_NUM79_OUT));
      NOR2_X1 XNOR_1_4_NUM79 (.ZN (XNOR_1_4_NUM79_OUT), .A1 (N320), .A2 (N352));
      NOR2_X1 XNOR_1_5_NUM79 (.ZN (N432), .A1 (XNOR_1_3_NUM79_OUT), .A2 (XNOR_1_4_NUM79_OUT));
      wire XNOR_1_1_NUM80_OUT, XNOR_1_2_NUM80_OUT, XNOR_1_3_NUM80_OUT, XNOR_1_4_NUM80_OUT;
      NOR2_X1 XNOR_1_1_NUM80 (.ZN (XNOR_1_1_NUM80_OUT), .A1 (N321), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM80 (.ZN (XNOR_1_2_NUM80_OUT), .A1 (GND), .A2 (N353));
      NOR2_X1 XNOR_1_3_NUM80 (.ZN (XNOR_1_3_NUM80_OUT), .A1 (XNOR_1_1_NUM80_OUT), .A2 (XNOR_1_2_NUM80_OUT));
      NOR2_X1 XNOR_1_4_NUM80 (.ZN (XNOR_1_4_NUM80_OUT), .A1 (N321), .A2 (N353));
      NOR2_X1 XNOR_1_5_NUM80 (.ZN (N445), .A1 (XNOR_1_3_NUM80_OUT), .A2 (XNOR_1_4_NUM80_OUT));
      NOR2_X1 XNOR_NUM81 (.ZN (N554), .A1 (N354), .A2 (GND));
      NOR2_X1 XNOR_NUM82 (.ZN (N555), .A1 (N367), .A2 (GND));
      NOR2_X1 XNOR_NUM83 (.ZN (N556), .A1 (N380), .A2 (GND));
      NOR2_X1 XNOR_NUM84 (.ZN (N557), .A1 (N354), .A2 (GND));
      NOR2_X1 XNOR_NUM85 (.ZN (N558), .A1 (N367), .A2 (GND));
      NOR2_X1 XNOR_NUM86 (.ZN (N559), .A1 (N393), .A2 (GND));
      NOR2_X1 XNOR_NUM87 (.ZN (N560), .A1 (N354), .A2 (GND));
      NOR2_X1 XNOR_NUM88 (.ZN (N561), .A1 (N380), .A2 (GND));
      NOR2_X1 XNOR_NUM89 (.ZN (N562), .A1 (N393), .A2 (GND));
      NOR2_X1 XNOR_NUM90 (.ZN (N563), .A1 (N367), .A2 (GND));
      NOR2_X1 XNOR_NUM91 (.ZN (N564), .A1 (N380), .A2 (GND));
      NOR2_X1 XNOR_NUM92 (.ZN (N565), .A1 (N393), .A2 (GND));
      NOR2_X1 XNOR_NUM93 (.ZN (N566), .A1 (N419), .A2 (GND));
      NOR2_X1 XNOR_NUM94 (.ZN (N567), .A1 (N445), .A2 (GND));
      NOR2_X1 XNOR_NUM95 (.ZN (N568), .A1 (N419), .A2 (GND));
      NOR2_X1 XNOR_NUM96 (.ZN (N569), .A1 (N432), .A2 (GND));
      NOR2_X1 XNOR_NUM97 (.ZN (N570), .A1 (N406), .A2 (GND));
      NOR2_X1 XNOR_NUM98 (.ZN (N571), .A1 (N445), .A2 (GND));
      NOR2_X1 XNOR_NUM99 (.ZN (N572), .A1 (N406), .A2 (GND));
      NOR2_X1 XNOR_NUM100 (.ZN (N573), .A1 (N432), .A2 (GND));
      NOR2_X1 XNOR_NUM101 (.ZN (N574), .A1 (N406), .A2 (GND));
      NOR2_X1 XNOR_NUM102 (.ZN (N575), .A1 (N419), .A2 (GND));
      NOR2_X1 XNOR_NUM103 (.ZN (N576), .A1 (N432), .A2 (GND));
      NOR2_X1 XNOR_NUM104 (.ZN (N577), .A1 (N406), .A2 (GND));
      NOR2_X1 XNOR_NUM105 (.ZN (N578), .A1 (N419), .A2 (GND));
      NOR2_X1 XNOR_NUM106 (.ZN (N579), .A1 (N445), .A2 (GND));
      NOR2_X1 XNOR_NUM107 (.ZN (N580), .A1 (N406), .A2 (GND));
      NOR2_X1 XNOR_NUM108 (.ZN (N581), .A1 (N432), .A2 (GND));
      NOR2_X1 XNOR_NUM109 (.ZN (N582), .A1 (N445), .A2 (GND));
      NOR2_X1 XNOR_NUM110 (.ZN (N583), .A1 (N419), .A2 (GND));
      NOR2_X1 XNOR_NUM111 (.ZN (N584), .A1 (N432), .A2 (GND));
      NOR2_X1 XNOR_NUM112 (.ZN (N585), .A1 (N445), .A2 (GND));
      NOR2_X1 XNOR_NUM113 (.ZN (N586), .A1 (N367), .A2 (GND));
      NOR2_X1 XNOR_NUM114 (.ZN (N587), .A1 (N393), .A2 (GND));
      NOR2_X1 XNOR_NUM115 (.ZN (N588), .A1 (N367), .A2 (GND));
      NOR2_X1 XNOR_NUM116 (.ZN (N589), .A1 (N380), .A2 (GND));
      NOR2_X1 XNOR_NUM117 (.ZN (N590), .A1 (N354), .A2 (GND));
      NOR2_X1 XNOR_NUM118 (.ZN (N591), .A1 (N393), .A2 (GND));
      NOR2_X1 XNOR_NUM119 (.ZN (N592), .A1 (N354), .A2 (GND));
      NOR2_X1 XNOR_NUM120 (.ZN (N593), .A1 (N380), .A2 (GND));
      wire XNOR_1_1_NUM121_OUT, XNOR_1_2_NUM121_OUT, XNOR_1_3_NUM121_OUT;
      NOR2_X1 XNOR_1_1_NUM121 (.ZN (XNOR_1_1_NUM121_OUT), .A1 (N554), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM121 (.ZN (XNOR_1_2_NUM121_OUT), .A1 (GND), .A2 (N555));
      NOR2_X1 XNOR_1_3_NUM121 (.ZN (XNOR_1_3_NUM121_OUT), .A1 (XNOR_1_1_NUM121_OUT), .A2 (XNOR_1_2_NUM121_OUT));

      wire XNOR_2_1_NUM121_OUT, XNOR_2_2_NUM121_OUT, XNOR_2_3_NUM121_OUT;
      NOR2_X1 XNOR_2_1_NUM121 (.ZN (XNOR_2_1_NUM121_OUT), .A1 (N556), .A2 (GND));
      NOR2_X1 XNOR_2_2_NUM121 (.ZN (XNOR_2_2_NUM121_OUT), .A1 (GND), .A2 (N393));
      NOR2_X1 XNOR_2_3_NUM121 (.ZN (XNOR_2_3_NUM121_OUT), .A1 (XNOR_2_1_NUM121_OUT), .A2 (XNOR_2_2_NUM121_OUT));

      wire XNOR_3_1_NUM121_OUT, XNOR_3_2_NUM121_OUT;
      NOR2_X1 XNOR_3_1_NUM121 (.ZN (XNOR_3_1_NUM121_OUT), .A1 (XNOR_1_3_NUM121_OUT), .A2 (GND));
      NOR2_X1 XNOR_3_2_NUM121 (.ZN (XNOR_3_2_NUM121_OUT), .A1 (GND), .A2 (XNOR_2_3_NUM121_OUT));
      NOR2_X1 XNOR_3_3_NUM121 (.ZN (N594), .A1 (XNOR_3_1_NUM121_OUT), .A2 (XNOR_3_2_NUM121_OUT));
      wire XNOR_1_1_NUM122_OUT, XNOR_1_2_NUM122_OUT, XNOR_1_3_NUM122_OUT;
      NOR2_X1 XNOR_1_1_NUM122 (.ZN (XNOR_1_1_NUM122_OUT), .A1 (N557), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM122 (.ZN (XNOR_1_2_NUM122_OUT), .A1 (GND), .A2 (N558));
      NOR2_X1 XNOR_1_3_NUM122 (.ZN (XNOR_1_3_NUM122_OUT), .A1 (XNOR_1_1_NUM122_OUT), .A2 (XNOR_1_2_NUM122_OUT));

      wire XNOR_2_1_NUM122_OUT, XNOR_2_2_NUM122_OUT, XNOR_2_3_NUM122_OUT;
      NOR2_X1 XNOR_2_1_NUM122 (.ZN (XNOR_2_1_NUM122_OUT), .A1 (N380), .A2 (GND));
      NOR2_X1 XNOR_2_2_NUM122 (.ZN (XNOR_2_2_NUM122_OUT), .A1 (GND), .A2 (N559));
      NOR2_X1 XNOR_2_3_NUM122 (.ZN (XNOR_2_3_NUM122_OUT), .A1 (XNOR_2_1_NUM122_OUT), .A2 (XNOR_2_2_NUM122_OUT));

      wire XNOR_3_1_NUM122_OUT, XNOR_3_2_NUM122_OUT;
      NOR2_X1 XNOR_3_1_NUM122 (.ZN (XNOR_3_1_NUM122_OUT), .A1 (XNOR_1_3_NUM122_OUT), .A2 (GND));
      NOR2_X1 XNOR_3_2_NUM122 (.ZN (XNOR_3_2_NUM122_OUT), .A1 (GND), .A2 (XNOR_2_3_NUM122_OUT));
      NOR2_X1 XNOR_3_3_NUM122 (.ZN (N595), .A1 (XNOR_3_1_NUM122_OUT), .A2 (XNOR_3_2_NUM122_OUT));
      wire XNOR_1_1_NUM123_OUT, XNOR_1_2_NUM123_OUT, XNOR_1_3_NUM123_OUT;
      NOR2_X1 XNOR_1_1_NUM123 (.ZN (XNOR_1_1_NUM123_OUT), .A1 (N560), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM123 (.ZN (XNOR_1_2_NUM123_OUT), .A1 (GND), .A2 (N367));
      NOR2_X1 XNOR_1_3_NUM123 (.ZN (XNOR_1_3_NUM123_OUT), .A1 (XNOR_1_1_NUM123_OUT), .A2 (XNOR_1_2_NUM123_OUT));

      wire XNOR_2_1_NUM123_OUT, XNOR_2_2_NUM123_OUT, XNOR_2_3_NUM123_OUT;
      NOR2_X1 XNOR_2_1_NUM123 (.ZN (XNOR_2_1_NUM123_OUT), .A1 (N561), .A2 (GND));
      NOR2_X1 XNOR_2_2_NUM123 (.ZN (XNOR_2_2_NUM123_OUT), .A1 (GND), .A2 (N562));
      NOR2_X1 XNOR_2_3_NUM123 (.ZN (XNOR_2_3_NUM123_OUT), .A1 (XNOR_2_1_NUM123_OUT), .A2 (XNOR_2_2_NUM123_OUT));

      wire XNOR_3_1_NUM123_OUT, XNOR_3_2_NUM123_OUT;
      NOR2_X1 XNOR_3_1_NUM123 (.ZN (XNOR_3_1_NUM123_OUT), .A1 (XNOR_1_3_NUM123_OUT), .A2 (GND));
      NOR2_X1 XNOR_3_2_NUM123 (.ZN (XNOR_3_2_NUM123_OUT), .A1 (GND), .A2 (XNOR_2_3_NUM123_OUT));
      NOR2_X1 XNOR_3_3_NUM123 (.ZN (N596), .A1 (XNOR_3_1_NUM123_OUT), .A2 (XNOR_3_2_NUM123_OUT));
      wire XNOR_1_1_NUM124_OUT, XNOR_1_2_NUM124_OUT, XNOR_1_3_NUM124_OUT;
      NOR2_X1 XNOR_1_1_NUM124 (.ZN (XNOR_1_1_NUM124_OUT), .A1 (N354), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM124 (.ZN (XNOR_1_2_NUM124_OUT), .A1 (GND), .A2 (N563));
      NOR2_X1 XNOR_1_3_NUM124 (.ZN (XNOR_1_3_NUM124_OUT), .A1 (XNOR_1_1_NUM124_OUT), .A2 (XNOR_1_2_NUM124_OUT));

      wire XNOR_2_1_NUM124_OUT, XNOR_2_2_NUM124_OUT, XNOR_2_3_NUM124_OUT;
      NOR2_X1 XNOR_2_1_NUM124 (.ZN (XNOR_2_1_NUM124_OUT), .A1 (N564), .A2 (GND));
      NOR2_X1 XNOR_2_2_NUM124 (.ZN (XNOR_2_2_NUM124_OUT), .A1 (GND), .A2 (N565));
      NOR2_X1 XNOR_2_3_NUM124 (.ZN (XNOR_2_3_NUM124_OUT), .A1 (XNOR_2_1_NUM124_OUT), .A2 (XNOR_2_2_NUM124_OUT));

      wire XNOR_3_1_NUM124_OUT, XNOR_3_2_NUM124_OUT;
      NOR2_X1 XNOR_3_1_NUM124 (.ZN (XNOR_3_1_NUM124_OUT), .A1 (XNOR_1_3_NUM124_OUT), .A2 (GND));
      NOR2_X1 XNOR_3_2_NUM124 (.ZN (XNOR_3_2_NUM124_OUT), .A1 (GND), .A2 (XNOR_2_3_NUM124_OUT));
      NOR2_X1 XNOR_3_3_NUM124 (.ZN (N597), .A1 (XNOR_3_1_NUM124_OUT), .A2 (XNOR_3_2_NUM124_OUT));
      wire XNOR_1_1_NUM125_OUT, XNOR_1_2_NUM125_OUT, XNOR_1_3_NUM125_OUT;
      NOR2_X1 XNOR_1_1_NUM125 (.ZN (XNOR_1_1_NUM125_OUT), .A1 (N574), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM125 (.ZN (XNOR_1_2_NUM125_OUT), .A1 (GND), .A2 (N575));
      NOR2_X1 XNOR_1_3_NUM125 (.ZN (XNOR_1_3_NUM125_OUT), .A1 (XNOR_1_1_NUM125_OUT), .A2 (XNOR_1_2_NUM125_OUT));

      wire XNOR_2_1_NUM125_OUT, XNOR_2_2_NUM125_OUT, XNOR_2_3_NUM125_OUT;
      NOR2_X1 XNOR_2_1_NUM125 (.ZN (XNOR_2_1_NUM125_OUT), .A1 (N576), .A2 (GND));
      NOR2_X1 XNOR_2_2_NUM125 (.ZN (XNOR_2_2_NUM125_OUT), .A1 (GND), .A2 (N445));
      NOR2_X1 XNOR_2_3_NUM125 (.ZN (XNOR_2_3_NUM125_OUT), .A1 (XNOR_2_1_NUM125_OUT), .A2 (XNOR_2_2_NUM125_OUT));

      wire XNOR_3_1_NUM125_OUT, XNOR_3_2_NUM125_OUT;
      NOR2_X1 XNOR_3_1_NUM125 (.ZN (XNOR_3_1_NUM125_OUT), .A1 (XNOR_1_3_NUM125_OUT), .A2 (GND));
      NOR2_X1 XNOR_3_2_NUM125 (.ZN (XNOR_3_2_NUM125_OUT), .A1 (GND), .A2 (XNOR_2_3_NUM125_OUT));
      NOR2_X1 XNOR_3_3_NUM125 (.ZN (N598), .A1 (XNOR_3_1_NUM125_OUT), .A2 (XNOR_3_2_NUM125_OUT));
      wire XNOR_1_1_NUM126_OUT, XNOR_1_2_NUM126_OUT, XNOR_1_3_NUM126_OUT;
      NOR2_X1 XNOR_1_1_NUM126 (.ZN (XNOR_1_1_NUM126_OUT), .A1 (N577), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM126 (.ZN (XNOR_1_2_NUM126_OUT), .A1 (GND), .A2 (N578));
      NOR2_X1 XNOR_1_3_NUM126 (.ZN (XNOR_1_3_NUM126_OUT), .A1 (XNOR_1_1_NUM126_OUT), .A2 (XNOR_1_2_NUM126_OUT));

      wire XNOR_2_1_NUM126_OUT, XNOR_2_2_NUM126_OUT, XNOR_2_3_NUM126_OUT;
      NOR2_X1 XNOR_2_1_NUM126 (.ZN (XNOR_2_1_NUM126_OUT), .A1 (N432), .A2 (GND));
      NOR2_X1 XNOR_2_2_NUM126 (.ZN (XNOR_2_2_NUM126_OUT), .A1 (GND), .A2 (N579));
      NOR2_X1 XNOR_2_3_NUM126 (.ZN (XNOR_2_3_NUM126_OUT), .A1 (XNOR_2_1_NUM126_OUT), .A2 (XNOR_2_2_NUM126_OUT));

      wire XNOR_3_1_NUM126_OUT, XNOR_3_2_NUM126_OUT;
      NOR2_X1 XNOR_3_1_NUM126 (.ZN (XNOR_3_1_NUM126_OUT), .A1 (XNOR_1_3_NUM126_OUT), .A2 (GND));
      NOR2_X1 XNOR_3_2_NUM126 (.ZN (XNOR_3_2_NUM126_OUT), .A1 (GND), .A2 (XNOR_2_3_NUM126_OUT));
      NOR2_X1 XNOR_3_3_NUM126 (.ZN (N599), .A1 (XNOR_3_1_NUM126_OUT), .A2 (XNOR_3_2_NUM126_OUT));
      wire XNOR_1_1_NUM127_OUT, XNOR_1_2_NUM127_OUT, XNOR_1_3_NUM127_OUT;
      NOR2_X1 XNOR_1_1_NUM127 (.ZN (XNOR_1_1_NUM127_OUT), .A1 (N580), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM127 (.ZN (XNOR_1_2_NUM127_OUT), .A1 (GND), .A2 (N419));
      NOR2_X1 XNOR_1_3_NUM127 (.ZN (XNOR_1_3_NUM127_OUT), .A1 (XNOR_1_1_NUM127_OUT), .A2 (XNOR_1_2_NUM127_OUT));

      wire XNOR_2_1_NUM127_OUT, XNOR_2_2_NUM127_OUT, XNOR_2_3_NUM127_OUT;
      NOR2_X1 XNOR_2_1_NUM127 (.ZN (XNOR_2_1_NUM127_OUT), .A1 (N581), .A2 (GND));
      NOR2_X1 XNOR_2_2_NUM127 (.ZN (XNOR_2_2_NUM127_OUT), .A1 (GND), .A2 (N582));
      NOR2_X1 XNOR_2_3_NUM127 (.ZN (XNOR_2_3_NUM127_OUT), .A1 (XNOR_2_1_NUM127_OUT), .A2 (XNOR_2_2_NUM127_OUT));

      wire XNOR_3_1_NUM127_OUT, XNOR_3_2_NUM127_OUT;
      NOR2_X1 XNOR_3_1_NUM127 (.ZN (XNOR_3_1_NUM127_OUT), .A1 (XNOR_1_3_NUM127_OUT), .A2 (GND));
      NOR2_X1 XNOR_3_2_NUM127 (.ZN (XNOR_3_2_NUM127_OUT), .A1 (GND), .A2 (XNOR_2_3_NUM127_OUT));
      NOR2_X1 XNOR_3_3_NUM127 (.ZN (N600), .A1 (XNOR_3_1_NUM127_OUT), .A2 (XNOR_3_2_NUM127_OUT));
      wire XNOR_1_1_NUM128_OUT, XNOR_1_2_NUM128_OUT, XNOR_1_3_NUM128_OUT;
      NOR2_X1 XNOR_1_1_NUM128 (.ZN (XNOR_1_1_NUM128_OUT), .A1 (N406), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM128 (.ZN (XNOR_1_2_NUM128_OUT), .A1 (GND), .A2 (N583));
      NOR2_X1 XNOR_1_3_NUM128 (.ZN (XNOR_1_3_NUM128_OUT), .A1 (XNOR_1_1_NUM128_OUT), .A2 (XNOR_1_2_NUM128_OUT));

      wire XNOR_2_1_NUM128_OUT, XNOR_2_2_NUM128_OUT, XNOR_2_3_NUM128_OUT;
      NOR2_X1 XNOR_2_1_NUM128 (.ZN (XNOR_2_1_NUM128_OUT), .A1 (N584), .A2 (GND));
      NOR2_X1 XNOR_2_2_NUM128 (.ZN (XNOR_2_2_NUM128_OUT), .A1 (GND), .A2 (N585));
      NOR2_X1 XNOR_2_3_NUM128 (.ZN (XNOR_2_3_NUM128_OUT), .A1 (XNOR_2_1_NUM128_OUT), .A2 (XNOR_2_2_NUM128_OUT));

      wire XNOR_3_1_NUM128_OUT, XNOR_3_2_NUM128_OUT;
      NOR2_X1 XNOR_3_1_NUM128 (.ZN (XNOR_3_1_NUM128_OUT), .A1 (XNOR_1_3_NUM128_OUT), .A2 (GND));
      NOR2_X1 XNOR_3_2_NUM128 (.ZN (XNOR_3_2_NUM128_OUT), .A1 (GND), .A2 (XNOR_2_3_NUM128_OUT));
      NOR2_X1 XNOR_3_3_NUM128 (.ZN (N601), .A1 (XNOR_3_1_NUM128_OUT), .A2 (XNOR_3_2_NUM128_OUT));
      wire XNOR_1_1_NUM129_OUT, XNOR_1_2_NUM129_OUT, XNOR_2_1_NUM129_OUT, XNOR_2_2_NUM129_OUT, XNOR_3_1_NUM129_OUT;
      NOR2_X1 XNOR_1_1_NUM129 (.ZN (XNOR_1_1_NUM129_OUT), .A1 (N594), .A2 (N595));
      NOR2_X1 XNOR_1_2_NUM129 (.ZN (XNOR_1_2_NUM129_OUT), .A1 (XNOR_1_1_NUM129_OUT), .A2 (GND));

      NOR2_X1 XNOR_2_1_NUM129 (.ZN (XNOR_2_1_NUM129_OUT), .A1 (N596), .A2 (N597));
      NOR2_X1 XNOR_2_2_NUM129 (.ZN (XNOR_2_2_NUM129_OUT), .A1 (XNOR_2_1_NUM129_OUT), .A2 (GND));

      NOR2_X1 XNOR_3_1_NUM129 (.ZN (XNOR_3_1_NUM129_OUT), .A1 (XNOR_1_2_NUM129_OUT), .A2 (XNOR_2_2_NUM129_OUT));
      NOR2_X1 XNOR_3_2_NUM129 (.ZN (N602), .A1 (XNOR_3_1_NUM129_OUT), .A2 (GND));
      wire XNOR_1_1_NUM130_OUT, XNOR_1_2_NUM130_OUT, XNOR_2_1_NUM130_OUT, XNOR_2_2_NUM130_OUT, XNOR_3_1_NUM130_OUT;
      NOR2_X1 XNOR_1_1_NUM130 (.ZN (XNOR_1_1_NUM130_OUT), .A1 (N598), .A2 (N599));
      NOR2_X1 XNOR_1_2_NUM130 (.ZN (XNOR_1_2_NUM130_OUT), .A1 (XNOR_1_1_NUM130_OUT), .A2 (GND));

      NOR2_X1 XNOR_2_1_NUM130 (.ZN (XNOR_2_1_NUM130_OUT), .A1 (N600), .A2 (N601));
      NOR2_X1 XNOR_2_2_NUM130 (.ZN (XNOR_2_2_NUM130_OUT), .A1 (XNOR_2_1_NUM130_OUT), .A2 (GND));

      NOR2_X1 XNOR_3_1_NUM130 (.ZN (XNOR_3_1_NUM130_OUT), .A1 (XNOR_1_2_NUM130_OUT), .A2 (XNOR_2_2_NUM130_OUT));
      NOR2_X1 XNOR_3_2_NUM130 (.ZN (N607), .A1 (XNOR_3_1_NUM130_OUT), .A2 (GND));
      wire XNOR_1_1_NUM131_OUT, XNOR_1_2_NUM131_OUT, XNOR_1_3_NUM131_OUT;
      NOR2_X1 XNOR_1_1_NUM131 (.ZN (XNOR_1_1_NUM131_OUT), .A1 (N406), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM131 (.ZN (XNOR_1_2_NUM131_OUT), .A1 (GND), .A2 (N566));
      NOR2_X1 XNOR_1_3_NUM131 (.ZN (XNOR_1_3_NUM131_OUT), .A1 (XNOR_1_1_NUM131_OUT), .A2 (XNOR_1_2_NUM131_OUT));

      wire XNOR_2_1_NUM131_OUT, XNOR_2_2_NUM131_OUT, XNOR_2_3_NUM131_OUT;
      NOR2_X1 XNOR_2_1_NUM131 (.ZN (XNOR_2_1_NUM131_OUT), .A1 (N432), .A2 (GND));
      NOR2_X1 XNOR_2_2_NUM131 (.ZN (XNOR_2_2_NUM131_OUT), .A1 (GND), .A2 (N567));
      NOR2_X1 XNOR_2_3_NUM131 (.ZN (XNOR_2_3_NUM131_OUT), .A1 (XNOR_2_1_NUM131_OUT), .A2 (XNOR_2_2_NUM131_OUT));

      wire XNOR_3_1_NUM131_OUT, XNOR_3_2_NUM131_OUT, XNOR_3_3_NUM131_OUT;
      NOR2_X1 XNOR_3_1_NUM131 (.ZN (XNOR_3_1_NUM131_OUT), .A1 (XNOR_1_3_NUM131_OUT), .A2 (GND));
      NOR2_X1 XNOR_3_2_NUM131 (.ZN (XNOR_3_2_NUM131_OUT), .A1 (GND), .A2 (XNOR_2_3_NUM131_OUT));
      NOR2_X1 XNOR_3_3_NUM131 (.ZN (XNOR_3_3_NUM131_OUT), .A1 (XNOR_3_1_NUM131_OUT), .A2 (XNOR_3_2_NUM131_OUT));

      wire XNOR_4_1_NUM131_OUT, XNOR_4_2_NUM131_OUT;
      NOR2_X1 XNOR_4_1_NUM131 (.ZN (XNOR_4_1_NUM131_OUT), .A1 (N602), .A2 (GND));
      NOR2_X1 XNOR_4_2_NUM131 (.ZN (XNOR_4_2_NUM131_OUT), .A1 (GND), .A2 (XNOR_3_3_NUM131_OUT));
      NOR2_X1 XNOR_4_3_NUM131 (.ZN (N620), .A1 (XNOR_4_1_NUM131_OUT), .A2 (XNOR_4_2_NUM131_OUT));
      wire XNOR_1_1_NUM132_OUT, XNOR_1_2_NUM132_OUT, XNOR_1_3_NUM132_OUT;
      NOR2_X1 XNOR_1_1_NUM132 (.ZN (XNOR_1_1_NUM132_OUT), .A1 (N406), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM132 (.ZN (XNOR_1_2_NUM132_OUT), .A1 (GND), .A2 (N568));
      NOR2_X1 XNOR_1_3_NUM132 (.ZN (XNOR_1_3_NUM132_OUT), .A1 (XNOR_1_1_NUM132_OUT), .A2 (XNOR_1_2_NUM132_OUT));

      wire XNOR_2_1_NUM132_OUT, XNOR_2_2_NUM132_OUT, XNOR_2_3_NUM132_OUT;
      NOR2_X1 XNOR_2_1_NUM132 (.ZN (XNOR_2_1_NUM132_OUT), .A1 (N569), .A2 (GND));
      NOR2_X1 XNOR_2_2_NUM132 (.ZN (XNOR_2_2_NUM132_OUT), .A1 (GND), .A2 (N445));
      NOR2_X1 XNOR_2_3_NUM132 (.ZN (XNOR_2_3_NUM132_OUT), .A1 (XNOR_2_1_NUM132_OUT), .A2 (XNOR_2_2_NUM132_OUT));

      wire XNOR_3_1_NUM132_OUT, XNOR_3_2_NUM132_OUT, XNOR_3_3_NUM132_OUT;
      NOR2_X1 XNOR_3_1_NUM132 (.ZN (XNOR_3_1_NUM132_OUT), .A1 (XNOR_1_3_NUM132_OUT), .A2 (GND));
      NOR2_X1 XNOR_3_2_NUM132 (.ZN (XNOR_3_2_NUM132_OUT), .A1 (GND), .A2 (XNOR_2_3_NUM132_OUT));
      NOR2_X1 XNOR_3_3_NUM132 (.ZN (XNOR_3_3_NUM132_OUT), .A1 (XNOR_3_1_NUM132_OUT), .A2 (XNOR_3_2_NUM132_OUT));

      wire XNOR_4_1_NUM132_OUT, XNOR_4_2_NUM132_OUT;
      NOR2_X1 XNOR_4_1_NUM132 (.ZN (XNOR_4_1_NUM132_OUT), .A1 (N602), .A2 (GND));
      NOR2_X1 XNOR_4_2_NUM132 (.ZN (XNOR_4_2_NUM132_OUT), .A1 (GND), .A2 (XNOR_3_3_NUM132_OUT));
      NOR2_X1 XNOR_4_3_NUM132 (.ZN (N625), .A1 (XNOR_4_1_NUM132_OUT), .A2 (XNOR_4_2_NUM132_OUT));
      wire XNOR_1_1_NUM133_OUT, XNOR_1_2_NUM133_OUT, XNOR_1_3_NUM133_OUT;
      NOR2_X1 XNOR_1_1_NUM133 (.ZN (XNOR_1_1_NUM133_OUT), .A1 (N570), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM133 (.ZN (XNOR_1_2_NUM133_OUT), .A1 (GND), .A2 (N419));
      NOR2_X1 XNOR_1_3_NUM133 (.ZN (XNOR_1_3_NUM133_OUT), .A1 (XNOR_1_1_NUM133_OUT), .A2 (XNOR_1_2_NUM133_OUT));

      wire XNOR_2_1_NUM133_OUT, XNOR_2_2_NUM133_OUT, XNOR_2_3_NUM133_OUT;
      NOR2_X1 XNOR_2_1_NUM133 (.ZN (XNOR_2_1_NUM133_OUT), .A1 (N432), .A2 (GND));
      NOR2_X1 XNOR_2_2_NUM133 (.ZN (XNOR_2_2_NUM133_OUT), .A1 (GND), .A2 (N571));
      NOR2_X1 XNOR_2_3_NUM133 (.ZN (XNOR_2_3_NUM133_OUT), .A1 (XNOR_2_1_NUM133_OUT), .A2 (XNOR_2_2_NUM133_OUT));

      wire XNOR_3_1_NUM133_OUT, XNOR_3_2_NUM133_OUT, XNOR_3_3_NUM133_OUT;
      NOR2_X1 XNOR_3_1_NUM133 (.ZN (XNOR_3_1_NUM133_OUT), .A1 (XNOR_1_3_NUM133_OUT), .A2 (GND));
      NOR2_X1 XNOR_3_2_NUM133 (.ZN (XNOR_3_2_NUM133_OUT), .A1 (GND), .A2 (XNOR_2_3_NUM133_OUT));
      NOR2_X1 XNOR_3_3_NUM133 (.ZN (XNOR_3_3_NUM133_OUT), .A1 (XNOR_3_1_NUM133_OUT), .A2 (XNOR_3_2_NUM133_OUT));

      wire XNOR_4_1_NUM133_OUT, XNOR_4_2_NUM133_OUT;
      NOR2_X1 XNOR_4_1_NUM133 (.ZN (XNOR_4_1_NUM133_OUT), .A1 (N602), .A2 (GND));
      NOR2_X1 XNOR_4_2_NUM133 (.ZN (XNOR_4_2_NUM133_OUT), .A1 (GND), .A2 (XNOR_3_3_NUM133_OUT));
      NOR2_X1 XNOR_4_3_NUM133 (.ZN (N630), .A1 (XNOR_4_1_NUM133_OUT), .A2 (XNOR_4_2_NUM133_OUT));
      wire XNOR_1_1_NUM134_OUT, XNOR_1_2_NUM134_OUT, XNOR_1_3_NUM134_OUT;
      NOR2_X1 XNOR_1_1_NUM134 (.ZN (XNOR_1_1_NUM134_OUT), .A1 (N572), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM134 (.ZN (XNOR_1_2_NUM134_OUT), .A1 (GND), .A2 (N419));
      NOR2_X1 XNOR_1_3_NUM134 (.ZN (XNOR_1_3_NUM134_OUT), .A1 (XNOR_1_1_NUM134_OUT), .A2 (XNOR_1_2_NUM134_OUT));

      wire XNOR_2_1_NUM134_OUT, XNOR_2_2_NUM134_OUT, XNOR_2_3_NUM134_OUT;
      NOR2_X1 XNOR_2_1_NUM134 (.ZN (XNOR_2_1_NUM134_OUT), .A1 (N573), .A2 (GND));
      NOR2_X1 XNOR_2_2_NUM134 (.ZN (XNOR_2_2_NUM134_OUT), .A1 (GND), .A2 (N445));
      NOR2_X1 XNOR_2_3_NUM134 (.ZN (XNOR_2_3_NUM134_OUT), .A1 (XNOR_2_1_NUM134_OUT), .A2 (XNOR_2_2_NUM134_OUT));

      wire XNOR_3_1_NUM134_OUT, XNOR_3_2_NUM134_OUT, XNOR_3_3_NUM134_OUT;
      NOR2_X1 XNOR_3_1_NUM134 (.ZN (XNOR_3_1_NUM134_OUT), .A1 (XNOR_1_3_NUM134_OUT), .A2 (GND));
      NOR2_X1 XNOR_3_2_NUM134 (.ZN (XNOR_3_2_NUM134_OUT), .A1 (GND), .A2 (XNOR_2_3_NUM134_OUT));
      NOR2_X1 XNOR_3_3_NUM134 (.ZN (XNOR_3_3_NUM134_OUT), .A1 (XNOR_3_1_NUM134_OUT), .A2 (XNOR_3_2_NUM134_OUT));

      wire XNOR_4_1_NUM134_OUT, XNOR_4_2_NUM134_OUT;
      NOR2_X1 XNOR_4_1_NUM134 (.ZN (XNOR_4_1_NUM134_OUT), .A1 (N602), .A2 (GND));
      NOR2_X1 XNOR_4_2_NUM134 (.ZN (XNOR_4_2_NUM134_OUT), .A1 (GND), .A2 (XNOR_3_3_NUM134_OUT));
      NOR2_X1 XNOR_4_3_NUM134 (.ZN (N635), .A1 (XNOR_4_1_NUM134_OUT), .A2 (XNOR_4_2_NUM134_OUT));
      wire XNOR_1_1_NUM135_OUT, XNOR_1_2_NUM135_OUT, XNOR_1_3_NUM135_OUT;
      NOR2_X1 XNOR_1_1_NUM135 (.ZN (XNOR_1_1_NUM135_OUT), .A1 (N354), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM135 (.ZN (XNOR_1_2_NUM135_OUT), .A1 (GND), .A2 (N586));
      NOR2_X1 XNOR_1_3_NUM135 (.ZN (XNOR_1_3_NUM135_OUT), .A1 (XNOR_1_1_NUM135_OUT), .A2 (XNOR_1_2_NUM135_OUT));

      wire XNOR_2_1_NUM135_OUT, XNOR_2_2_NUM135_OUT, XNOR_2_3_NUM135_OUT;
      NOR2_X1 XNOR_2_1_NUM135 (.ZN (XNOR_2_1_NUM135_OUT), .A1 (N380), .A2 (GND));
      NOR2_X1 XNOR_2_2_NUM135 (.ZN (XNOR_2_2_NUM135_OUT), .A1 (GND), .A2 (N587));
      NOR2_X1 XNOR_2_3_NUM135 (.ZN (XNOR_2_3_NUM135_OUT), .A1 (XNOR_2_1_NUM135_OUT), .A2 (XNOR_2_2_NUM135_OUT));

      wire XNOR_3_1_NUM135_OUT, XNOR_3_2_NUM135_OUT, XNOR_3_3_NUM135_OUT;
      NOR2_X1 XNOR_3_1_NUM135 (.ZN (XNOR_3_1_NUM135_OUT), .A1 (XNOR_1_3_NUM135_OUT), .A2 (GND));
      NOR2_X1 XNOR_3_2_NUM135 (.ZN (XNOR_3_2_NUM135_OUT), .A1 (GND), .A2 (XNOR_2_3_NUM135_OUT));
      NOR2_X1 XNOR_3_3_NUM135 (.ZN (XNOR_3_3_NUM135_OUT), .A1 (XNOR_3_1_NUM135_OUT), .A2 (XNOR_3_2_NUM135_OUT));

      wire XNOR_4_1_NUM135_OUT, XNOR_4_2_NUM135_OUT;
      NOR2_X1 XNOR_4_1_NUM135 (.ZN (XNOR_4_1_NUM135_OUT), .A1 (N607), .A2 (GND));
      NOR2_X1 XNOR_4_2_NUM135 (.ZN (XNOR_4_2_NUM135_OUT), .A1 (GND), .A2 (XNOR_3_3_NUM135_OUT));
      NOR2_X1 XNOR_4_3_NUM135 (.ZN (N640), .A1 (XNOR_4_1_NUM135_OUT), .A2 (XNOR_4_2_NUM135_OUT));
      wire XNOR_1_1_NUM136_OUT, XNOR_1_2_NUM136_OUT, XNOR_1_3_NUM136_OUT;
      NOR2_X1 XNOR_1_1_NUM136 (.ZN (XNOR_1_1_NUM136_OUT), .A1 (N354), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM136 (.ZN (XNOR_1_2_NUM136_OUT), .A1 (GND), .A2 (N588));
      NOR2_X1 XNOR_1_3_NUM136 (.ZN (XNOR_1_3_NUM136_OUT), .A1 (XNOR_1_1_NUM136_OUT), .A2 (XNOR_1_2_NUM136_OUT));

      wire XNOR_2_1_NUM136_OUT, XNOR_2_2_NUM136_OUT, XNOR_2_3_NUM136_OUT;
      NOR2_X1 XNOR_2_1_NUM136 (.ZN (XNOR_2_1_NUM136_OUT), .A1 (N589), .A2 (GND));
      NOR2_X1 XNOR_2_2_NUM136 (.ZN (XNOR_2_2_NUM136_OUT), .A1 (GND), .A2 (N393));
      NOR2_X1 XNOR_2_3_NUM136 (.ZN (XNOR_2_3_NUM136_OUT), .A1 (XNOR_2_1_NUM136_OUT), .A2 (XNOR_2_2_NUM136_OUT));

      wire XNOR_3_1_NUM136_OUT, XNOR_3_2_NUM136_OUT, XNOR_3_3_NUM136_OUT;
      NOR2_X1 XNOR_3_1_NUM136 (.ZN (XNOR_3_1_NUM136_OUT), .A1 (XNOR_1_3_NUM136_OUT), .A2 (GND));
      NOR2_X1 XNOR_3_2_NUM136 (.ZN (XNOR_3_2_NUM136_OUT), .A1 (GND), .A2 (XNOR_2_3_NUM136_OUT));
      NOR2_X1 XNOR_3_3_NUM136 (.ZN (XNOR_3_3_NUM136_OUT), .A1 (XNOR_3_1_NUM136_OUT), .A2 (XNOR_3_2_NUM136_OUT));

      wire XNOR_4_1_NUM136_OUT, XNOR_4_2_NUM136_OUT;
      NOR2_X1 XNOR_4_1_NUM136 (.ZN (XNOR_4_1_NUM136_OUT), .A1 (N607), .A2 (GND));
      NOR2_X1 XNOR_4_2_NUM136 (.ZN (XNOR_4_2_NUM136_OUT), .A1 (GND), .A2 (XNOR_3_3_NUM136_OUT));
      NOR2_X1 XNOR_4_3_NUM136 (.ZN (N645), .A1 (XNOR_4_1_NUM136_OUT), .A2 (XNOR_4_2_NUM136_OUT));
      wire XNOR_1_1_NUM137_OUT, XNOR_1_2_NUM137_OUT, XNOR_1_3_NUM137_OUT;
      NOR2_X1 XNOR_1_1_NUM137 (.ZN (XNOR_1_1_NUM137_OUT), .A1 (N590), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM137 (.ZN (XNOR_1_2_NUM137_OUT), .A1 (GND), .A2 (N367));
      NOR2_X1 XNOR_1_3_NUM137 (.ZN (XNOR_1_3_NUM137_OUT), .A1 (XNOR_1_1_NUM137_OUT), .A2 (XNOR_1_2_NUM137_OUT));

      wire XNOR_2_1_NUM137_OUT, XNOR_2_2_NUM137_OUT, XNOR_2_3_NUM137_OUT;
      NOR2_X1 XNOR_2_1_NUM137 (.ZN (XNOR_2_1_NUM137_OUT), .A1 (N380), .A2 (GND));
      NOR2_X1 XNOR_2_2_NUM137 (.ZN (XNOR_2_2_NUM137_OUT), .A1 (GND), .A2 (N591));
      NOR2_X1 XNOR_2_3_NUM137 (.ZN (XNOR_2_3_NUM137_OUT), .A1 (XNOR_2_1_NUM137_OUT), .A2 (XNOR_2_2_NUM137_OUT));

      wire XNOR_3_1_NUM137_OUT, XNOR_3_2_NUM137_OUT, XNOR_3_3_NUM137_OUT;
      NOR2_X1 XNOR_3_1_NUM137 (.ZN (XNOR_3_1_NUM137_OUT), .A1 (XNOR_1_3_NUM137_OUT), .A2 (GND));
      NOR2_X1 XNOR_3_2_NUM137 (.ZN (XNOR_3_2_NUM137_OUT), .A1 (GND), .A2 (XNOR_2_3_NUM137_OUT));
      NOR2_X1 XNOR_3_3_NUM137 (.ZN (XNOR_3_3_NUM137_OUT), .A1 (XNOR_3_1_NUM137_OUT), .A2 (XNOR_3_2_NUM137_OUT));

      wire XNOR_4_1_NUM137_OUT, XNOR_4_2_NUM137_OUT;
      NOR2_X1 XNOR_4_1_NUM137 (.ZN (XNOR_4_1_NUM137_OUT), .A1 (N607), .A2 (GND));
      NOR2_X1 XNOR_4_2_NUM137 (.ZN (XNOR_4_2_NUM137_OUT), .A1 (GND), .A2 (XNOR_3_3_NUM137_OUT));
      NOR2_X1 XNOR_4_3_NUM137 (.ZN (N650), .A1 (XNOR_4_1_NUM137_OUT), .A2 (XNOR_4_2_NUM137_OUT));
      wire XNOR_1_1_NUM138_OUT, XNOR_1_2_NUM138_OUT, XNOR_1_3_NUM138_OUT;
      NOR2_X1 XNOR_1_1_NUM138 (.ZN (XNOR_1_1_NUM138_OUT), .A1 (N592), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM138 (.ZN (XNOR_1_2_NUM138_OUT), .A1 (GND), .A2 (N367));
      NOR2_X1 XNOR_1_3_NUM138 (.ZN (XNOR_1_3_NUM138_OUT), .A1 (XNOR_1_1_NUM138_OUT), .A2 (XNOR_1_2_NUM138_OUT));

      wire XNOR_2_1_NUM138_OUT, XNOR_2_2_NUM138_OUT, XNOR_2_3_NUM138_OUT;
      NOR2_X1 XNOR_2_1_NUM138 (.ZN (XNOR_2_1_NUM138_OUT), .A1 (N593), .A2 (GND));
      NOR2_X1 XNOR_2_2_NUM138 (.ZN (XNOR_2_2_NUM138_OUT), .A1 (GND), .A2 (N393));
      NOR2_X1 XNOR_2_3_NUM138 (.ZN (XNOR_2_3_NUM138_OUT), .A1 (XNOR_2_1_NUM138_OUT), .A2 (XNOR_2_2_NUM138_OUT));

      wire XNOR_3_1_NUM138_OUT, XNOR_3_2_NUM138_OUT, XNOR_3_3_NUM138_OUT;
      NOR2_X1 XNOR_3_1_NUM138 (.ZN (XNOR_3_1_NUM138_OUT), .A1 (XNOR_1_3_NUM138_OUT), .A2 (GND));
      NOR2_X1 XNOR_3_2_NUM138 (.ZN (XNOR_3_2_NUM138_OUT), .A1 (GND), .A2 (XNOR_2_3_NUM138_OUT));
      NOR2_X1 XNOR_3_3_NUM138 (.ZN (XNOR_3_3_NUM138_OUT), .A1 (XNOR_3_1_NUM138_OUT), .A2 (XNOR_3_2_NUM138_OUT));

      wire XNOR_4_1_NUM138_OUT, XNOR_4_2_NUM138_OUT;
      NOR2_X1 XNOR_4_1_NUM138 (.ZN (XNOR_4_1_NUM138_OUT), .A1 (N607), .A2 (GND));
      NOR2_X1 XNOR_4_2_NUM138 (.ZN (XNOR_4_2_NUM138_OUT), .A1 (GND), .A2 (XNOR_3_3_NUM138_OUT));
      NOR2_X1 XNOR_4_3_NUM138 (.ZN (N655), .A1 (XNOR_4_1_NUM138_OUT), .A2 (XNOR_4_2_NUM138_OUT));
      wire XNOR_1_1_NUM139_OUT, XNOR_1_2_NUM139_OUT;
      NOR2_X1 XNOR_1_1_NUM139 (.ZN (XNOR_1_1_NUM139_OUT), .A1 (N354), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM139 (.ZN (XNOR_1_2_NUM139_OUT), .A1 (GND), .A2 (N620));
      NOR2_X1 XNOR_1_3_NUM139 (.ZN (N692), .A1 (XNOR_1_1_NUM139_OUT), .A2 (XNOR_1_2_NUM139_OUT));
      wire XNOR_1_1_NUM140_OUT, XNOR_1_2_NUM140_OUT;
      NOR2_X1 XNOR_1_1_NUM140 (.ZN (XNOR_1_1_NUM140_OUT), .A1 (N367), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM140 (.ZN (XNOR_1_2_NUM140_OUT), .A1 (GND), .A2 (N620));
      NOR2_X1 XNOR_1_3_NUM140 (.ZN (N693), .A1 (XNOR_1_1_NUM140_OUT), .A2 (XNOR_1_2_NUM140_OUT));
      wire XNOR_1_1_NUM141_OUT, XNOR_1_2_NUM141_OUT;
      NOR2_X1 XNOR_1_1_NUM141 (.ZN (XNOR_1_1_NUM141_OUT), .A1 (N380), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM141 (.ZN (XNOR_1_2_NUM141_OUT), .A1 (GND), .A2 (N620));
      NOR2_X1 XNOR_1_3_NUM141 (.ZN (N694), .A1 (XNOR_1_1_NUM141_OUT), .A2 (XNOR_1_2_NUM141_OUT));
      wire XNOR_1_1_NUM142_OUT, XNOR_1_2_NUM142_OUT;
      NOR2_X1 XNOR_1_1_NUM142 (.ZN (XNOR_1_1_NUM142_OUT), .A1 (N393), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM142 (.ZN (XNOR_1_2_NUM142_OUT), .A1 (GND), .A2 (N620));
      NOR2_X1 XNOR_1_3_NUM142 (.ZN (N695), .A1 (XNOR_1_1_NUM142_OUT), .A2 (XNOR_1_2_NUM142_OUT));
      wire XNOR_1_1_NUM143_OUT, XNOR_1_2_NUM143_OUT;
      NOR2_X1 XNOR_1_1_NUM143 (.ZN (XNOR_1_1_NUM143_OUT), .A1 (N354), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM143 (.ZN (XNOR_1_2_NUM143_OUT), .A1 (GND), .A2 (N625));
      NOR2_X1 XNOR_1_3_NUM143 (.ZN (N696), .A1 (XNOR_1_1_NUM143_OUT), .A2 (XNOR_1_2_NUM143_OUT));
      wire XNOR_1_1_NUM144_OUT, XNOR_1_2_NUM144_OUT;
      NOR2_X1 XNOR_1_1_NUM144 (.ZN (XNOR_1_1_NUM144_OUT), .A1 (N367), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM144 (.ZN (XNOR_1_2_NUM144_OUT), .A1 (GND), .A2 (N625));
      NOR2_X1 XNOR_1_3_NUM144 (.ZN (N697), .A1 (XNOR_1_1_NUM144_OUT), .A2 (XNOR_1_2_NUM144_OUT));
      wire XNOR_1_1_NUM145_OUT, XNOR_1_2_NUM145_OUT;
      NOR2_X1 XNOR_1_1_NUM145 (.ZN (XNOR_1_1_NUM145_OUT), .A1 (N380), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM145 (.ZN (XNOR_1_2_NUM145_OUT), .A1 (GND), .A2 (N625));
      NOR2_X1 XNOR_1_3_NUM145 (.ZN (N698), .A1 (XNOR_1_1_NUM145_OUT), .A2 (XNOR_1_2_NUM145_OUT));
      wire XNOR_1_1_NUM146_OUT, XNOR_1_2_NUM146_OUT;
      NOR2_X1 XNOR_1_1_NUM146 (.ZN (XNOR_1_1_NUM146_OUT), .A1 (N393), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM146 (.ZN (XNOR_1_2_NUM146_OUT), .A1 (GND), .A2 (N625));
      NOR2_X1 XNOR_1_3_NUM146 (.ZN (N699), .A1 (XNOR_1_1_NUM146_OUT), .A2 (XNOR_1_2_NUM146_OUT));
      wire XNOR_1_1_NUM147_OUT, XNOR_1_2_NUM147_OUT;
      NOR2_X1 XNOR_1_1_NUM147 (.ZN (XNOR_1_1_NUM147_OUT), .A1 (N354), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM147 (.ZN (XNOR_1_2_NUM147_OUT), .A1 (GND), .A2 (N630));
      NOR2_X1 XNOR_1_3_NUM147 (.ZN (N700), .A1 (XNOR_1_1_NUM147_OUT), .A2 (XNOR_1_2_NUM147_OUT));
      wire XNOR_1_1_NUM148_OUT, XNOR_1_2_NUM148_OUT;
      NOR2_X1 XNOR_1_1_NUM148 (.ZN (XNOR_1_1_NUM148_OUT), .A1 (N367), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM148 (.ZN (XNOR_1_2_NUM148_OUT), .A1 (GND), .A2 (N630));
      NOR2_X1 XNOR_1_3_NUM148 (.ZN (N701), .A1 (XNOR_1_1_NUM148_OUT), .A2 (XNOR_1_2_NUM148_OUT));
      wire XNOR_1_1_NUM149_OUT, XNOR_1_2_NUM149_OUT;
      NOR2_X1 XNOR_1_1_NUM149 (.ZN (XNOR_1_1_NUM149_OUT), .A1 (N380), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM149 (.ZN (XNOR_1_2_NUM149_OUT), .A1 (GND), .A2 (N630));
      NOR2_X1 XNOR_1_3_NUM149 (.ZN (N702), .A1 (XNOR_1_1_NUM149_OUT), .A2 (XNOR_1_2_NUM149_OUT));
      wire XNOR_1_1_NUM150_OUT, XNOR_1_2_NUM150_OUT;
      NOR2_X1 XNOR_1_1_NUM150 (.ZN (XNOR_1_1_NUM150_OUT), .A1 (N393), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM150 (.ZN (XNOR_1_2_NUM150_OUT), .A1 (GND), .A2 (N630));
      NOR2_X1 XNOR_1_3_NUM150 (.ZN (N703), .A1 (XNOR_1_1_NUM150_OUT), .A2 (XNOR_1_2_NUM150_OUT));
      wire XNOR_1_1_NUM151_OUT, XNOR_1_2_NUM151_OUT;
      NOR2_X1 XNOR_1_1_NUM151 (.ZN (XNOR_1_1_NUM151_OUT), .A1 (N354), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM151 (.ZN (XNOR_1_2_NUM151_OUT), .A1 (GND), .A2 (N635));
      NOR2_X1 XNOR_1_3_NUM151 (.ZN (N704), .A1 (XNOR_1_1_NUM151_OUT), .A2 (XNOR_1_2_NUM151_OUT));
      wire XNOR_1_1_NUM152_OUT, XNOR_1_2_NUM152_OUT;
      NOR2_X1 XNOR_1_1_NUM152 (.ZN (XNOR_1_1_NUM152_OUT), .A1 (N367), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM152 (.ZN (XNOR_1_2_NUM152_OUT), .A1 (GND), .A2 (N635));
      NOR2_X1 XNOR_1_3_NUM152 (.ZN (N705), .A1 (XNOR_1_1_NUM152_OUT), .A2 (XNOR_1_2_NUM152_OUT));
      wire XNOR_1_1_NUM153_OUT, XNOR_1_2_NUM153_OUT;
      NOR2_X1 XNOR_1_1_NUM153 (.ZN (XNOR_1_1_NUM153_OUT), .A1 (N380), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM153 (.ZN (XNOR_1_2_NUM153_OUT), .A1 (GND), .A2 (N635));
      NOR2_X1 XNOR_1_3_NUM153 (.ZN (N706), .A1 (XNOR_1_1_NUM153_OUT), .A2 (XNOR_1_2_NUM153_OUT));
      wire XNOR_1_1_NUM154_OUT, XNOR_1_2_NUM154_OUT;
      NOR2_X1 XNOR_1_1_NUM154 (.ZN (XNOR_1_1_NUM154_OUT), .A1 (N393), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM154 (.ZN (XNOR_1_2_NUM154_OUT), .A1 (GND), .A2 (N635));
      NOR2_X1 XNOR_1_3_NUM154 (.ZN (N707), .A1 (XNOR_1_1_NUM154_OUT), .A2 (XNOR_1_2_NUM154_OUT));
      wire XNOR_1_1_NUM155_OUT, XNOR_1_2_NUM155_OUT;
      NOR2_X1 XNOR_1_1_NUM155 (.ZN (XNOR_1_1_NUM155_OUT), .A1 (N406), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM155 (.ZN (XNOR_1_2_NUM155_OUT), .A1 (GND), .A2 (N640));
      NOR2_X1 XNOR_1_3_NUM155 (.ZN (N708), .A1 (XNOR_1_1_NUM155_OUT), .A2 (XNOR_1_2_NUM155_OUT));
      wire XNOR_1_1_NUM156_OUT, XNOR_1_2_NUM156_OUT;
      NOR2_X1 XNOR_1_1_NUM156 (.ZN (XNOR_1_1_NUM156_OUT), .A1 (N419), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM156 (.ZN (XNOR_1_2_NUM156_OUT), .A1 (GND), .A2 (N640));
      NOR2_X1 XNOR_1_3_NUM156 (.ZN (N709), .A1 (XNOR_1_1_NUM156_OUT), .A2 (XNOR_1_2_NUM156_OUT));
      wire XNOR_1_1_NUM157_OUT, XNOR_1_2_NUM157_OUT;
      NOR2_X1 XNOR_1_1_NUM157 (.ZN (XNOR_1_1_NUM157_OUT), .A1 (N432), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM157 (.ZN (XNOR_1_2_NUM157_OUT), .A1 (GND), .A2 (N640));
      NOR2_X1 XNOR_1_3_NUM157 (.ZN (N710), .A1 (XNOR_1_1_NUM157_OUT), .A2 (XNOR_1_2_NUM157_OUT));
      wire XNOR_1_1_NUM158_OUT, XNOR_1_2_NUM158_OUT;
      NOR2_X1 XNOR_1_1_NUM158 (.ZN (XNOR_1_1_NUM158_OUT), .A1 (N445), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM158 (.ZN (XNOR_1_2_NUM158_OUT), .A1 (GND), .A2 (N640));
      NOR2_X1 XNOR_1_3_NUM158 (.ZN (N711), .A1 (XNOR_1_1_NUM158_OUT), .A2 (XNOR_1_2_NUM158_OUT));
      wire XNOR_1_1_NUM159_OUT, XNOR_1_2_NUM159_OUT;
      NOR2_X1 XNOR_1_1_NUM159 (.ZN (XNOR_1_1_NUM159_OUT), .A1 (N406), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM159 (.ZN (XNOR_1_2_NUM159_OUT), .A1 (GND), .A2 (N645));
      NOR2_X1 XNOR_1_3_NUM159 (.ZN (N712), .A1 (XNOR_1_1_NUM159_OUT), .A2 (XNOR_1_2_NUM159_OUT));
      wire XNOR_1_1_NUM160_OUT, XNOR_1_2_NUM160_OUT;
      NOR2_X1 XNOR_1_1_NUM160 (.ZN (XNOR_1_1_NUM160_OUT), .A1 (N419), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM160 (.ZN (XNOR_1_2_NUM160_OUT), .A1 (GND), .A2 (N645));
      NOR2_X1 XNOR_1_3_NUM160 (.ZN (N713), .A1 (XNOR_1_1_NUM160_OUT), .A2 (XNOR_1_2_NUM160_OUT));
      wire XNOR_1_1_NUM161_OUT, XNOR_1_2_NUM161_OUT;
      NOR2_X1 XNOR_1_1_NUM161 (.ZN (XNOR_1_1_NUM161_OUT), .A1 (N432), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM161 (.ZN (XNOR_1_2_NUM161_OUT), .A1 (GND), .A2 (N645));
      NOR2_X1 XNOR_1_3_NUM161 (.ZN (N714), .A1 (XNOR_1_1_NUM161_OUT), .A2 (XNOR_1_2_NUM161_OUT));
      wire XNOR_1_1_NUM162_OUT, XNOR_1_2_NUM162_OUT;
      NOR2_X1 XNOR_1_1_NUM162 (.ZN (XNOR_1_1_NUM162_OUT), .A1 (N445), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM162 (.ZN (XNOR_1_2_NUM162_OUT), .A1 (GND), .A2 (N645));
      NOR2_X1 XNOR_1_3_NUM162 (.ZN (N715), .A1 (XNOR_1_1_NUM162_OUT), .A2 (XNOR_1_2_NUM162_OUT));
      wire XNOR_1_1_NUM163_OUT, XNOR_1_2_NUM163_OUT;
      NOR2_X1 XNOR_1_1_NUM163 (.ZN (XNOR_1_1_NUM163_OUT), .A1 (N406), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM163 (.ZN (XNOR_1_2_NUM163_OUT), .A1 (GND), .A2 (N650));
      NOR2_X1 XNOR_1_3_NUM163 (.ZN (N716), .A1 (XNOR_1_1_NUM163_OUT), .A2 (XNOR_1_2_NUM163_OUT));
      wire XNOR_1_1_NUM164_OUT, XNOR_1_2_NUM164_OUT;
      NOR2_X1 XNOR_1_1_NUM164 (.ZN (XNOR_1_1_NUM164_OUT), .A1 (N419), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM164 (.ZN (XNOR_1_2_NUM164_OUT), .A1 (GND), .A2 (N650));
      NOR2_X1 XNOR_1_3_NUM164 (.ZN (N717), .A1 (XNOR_1_1_NUM164_OUT), .A2 (XNOR_1_2_NUM164_OUT));
      wire XNOR_1_1_NUM165_OUT, XNOR_1_2_NUM165_OUT;
      NOR2_X1 XNOR_1_1_NUM165 (.ZN (XNOR_1_1_NUM165_OUT), .A1 (N432), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM165 (.ZN (XNOR_1_2_NUM165_OUT), .A1 (GND), .A2 (N650));
      NOR2_X1 XNOR_1_3_NUM165 (.ZN (N718), .A1 (XNOR_1_1_NUM165_OUT), .A2 (XNOR_1_2_NUM165_OUT));
      wire XNOR_1_1_NUM166_OUT, XNOR_1_2_NUM166_OUT;
      NOR2_X1 XNOR_1_1_NUM166 (.ZN (XNOR_1_1_NUM166_OUT), .A1 (N445), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM166 (.ZN (XNOR_1_2_NUM166_OUT), .A1 (GND), .A2 (N650));
      NOR2_X1 XNOR_1_3_NUM166 (.ZN (N719), .A1 (XNOR_1_1_NUM166_OUT), .A2 (XNOR_1_2_NUM166_OUT));
      wire XNOR_1_1_NUM167_OUT, XNOR_1_2_NUM167_OUT;
      NOR2_X1 XNOR_1_1_NUM167 (.ZN (XNOR_1_1_NUM167_OUT), .A1 (N406), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM167 (.ZN (XNOR_1_2_NUM167_OUT), .A1 (GND), .A2 (N655));
      NOR2_X1 XNOR_1_3_NUM167 (.ZN (N720), .A1 (XNOR_1_1_NUM167_OUT), .A2 (XNOR_1_2_NUM167_OUT));
      wire XNOR_1_1_NUM168_OUT, XNOR_1_2_NUM168_OUT;
      NOR2_X1 XNOR_1_1_NUM168 (.ZN (XNOR_1_1_NUM168_OUT), .A1 (N419), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM168 (.ZN (XNOR_1_2_NUM168_OUT), .A1 (GND), .A2 (N655));
      NOR2_X1 XNOR_1_3_NUM168 (.ZN (N721), .A1 (XNOR_1_1_NUM168_OUT), .A2 (XNOR_1_2_NUM168_OUT));
      wire XNOR_1_1_NUM169_OUT, XNOR_1_2_NUM169_OUT;
      NOR2_X1 XNOR_1_1_NUM169 (.ZN (XNOR_1_1_NUM169_OUT), .A1 (N432), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM169 (.ZN (XNOR_1_2_NUM169_OUT), .A1 (GND), .A2 (N655));
      NOR2_X1 XNOR_1_3_NUM169 (.ZN (N722), .A1 (XNOR_1_1_NUM169_OUT), .A2 (XNOR_1_2_NUM169_OUT));
      wire XNOR_1_1_NUM170_OUT, XNOR_1_2_NUM170_OUT;
      NOR2_X1 XNOR_1_1_NUM170 (.ZN (XNOR_1_1_NUM170_OUT), .A1 (N445), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM170 (.ZN (XNOR_1_2_NUM170_OUT), .A1 (GND), .A2 (N655));
      NOR2_X1 XNOR_1_3_NUM170 (.ZN (N723), .A1 (XNOR_1_1_NUM170_OUT), .A2 (XNOR_1_2_NUM170_OUT));
      wire XNOR_1_1_NUM171_OUT, XNOR_1_2_NUM171_OUT, XNOR_1_3_NUM171_OUT, XNOR_1_4_NUM171_OUT;
      NOR2_X1 XNOR_1_1_NUM171 (.ZN (XNOR_1_1_NUM171_OUT), .A1 (N1), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM171 (.ZN (XNOR_1_2_NUM171_OUT), .A1 (GND), .A2 (N692));
      NOR2_X1 XNOR_1_3_NUM171 (.ZN (XNOR_1_3_NUM171_OUT), .A1 (XNOR_1_1_NUM171_OUT), .A2 (XNOR_1_2_NUM171_OUT));
      NOR2_X1 XNOR_1_4_NUM171 (.ZN (XNOR_1_4_NUM171_OUT), .A1 (N1), .A2 (N692));
      NOR2_X1 XNOR_1_5_NUM171 (.ZN (N724), .A1 (XNOR_1_3_NUM171_OUT), .A2 (XNOR_1_4_NUM171_OUT));
      wire XNOR_1_1_NUM172_OUT, XNOR_1_2_NUM172_OUT, XNOR_1_3_NUM172_OUT, XNOR_1_4_NUM172_OUT;
      NOR2_X1 XNOR_1_1_NUM172 (.ZN (XNOR_1_1_NUM172_OUT), .A1 (N5), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM172 (.ZN (XNOR_1_2_NUM172_OUT), .A1 (GND), .A2 (N693));
      NOR2_X1 XNOR_1_3_NUM172 (.ZN (XNOR_1_3_NUM172_OUT), .A1 (XNOR_1_1_NUM172_OUT), .A2 (XNOR_1_2_NUM172_OUT));
      NOR2_X1 XNOR_1_4_NUM172 (.ZN (XNOR_1_4_NUM172_OUT), .A1 (N5), .A2 (N693));
      NOR2_X1 XNOR_1_5_NUM172 (.ZN (N725), .A1 (XNOR_1_3_NUM172_OUT), .A2 (XNOR_1_4_NUM172_OUT));
      wire XNOR_1_1_NUM173_OUT, XNOR_1_2_NUM173_OUT, XNOR_1_3_NUM173_OUT, XNOR_1_4_NUM173_OUT;
      NOR2_X1 XNOR_1_1_NUM173 (.ZN (XNOR_1_1_NUM173_OUT), .A1 (N9), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM173 (.ZN (XNOR_1_2_NUM173_OUT), .A1 (GND), .A2 (N694));
      NOR2_X1 XNOR_1_3_NUM173 (.ZN (XNOR_1_3_NUM173_OUT), .A1 (XNOR_1_1_NUM173_OUT), .A2 (XNOR_1_2_NUM173_OUT));
      NOR2_X1 XNOR_1_4_NUM173 (.ZN (XNOR_1_4_NUM173_OUT), .A1 (N9), .A2 (N694));
      NOR2_X1 XNOR_1_5_NUM173 (.ZN (N726), .A1 (XNOR_1_3_NUM173_OUT), .A2 (XNOR_1_4_NUM173_OUT));
      wire XNOR_1_1_NUM174_OUT, XNOR_1_2_NUM174_OUT, XNOR_1_3_NUM174_OUT, XNOR_1_4_NUM174_OUT;
      NOR2_X1 XNOR_1_1_NUM174 (.ZN (XNOR_1_1_NUM174_OUT), .A1 (N13), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM174 (.ZN (XNOR_1_2_NUM174_OUT), .A1 (GND), .A2 (N695));
      NOR2_X1 XNOR_1_3_NUM174 (.ZN (XNOR_1_3_NUM174_OUT), .A1 (XNOR_1_1_NUM174_OUT), .A2 (XNOR_1_2_NUM174_OUT));
      NOR2_X1 XNOR_1_4_NUM174 (.ZN (XNOR_1_4_NUM174_OUT), .A1 (N13), .A2 (N695));
      NOR2_X1 XNOR_1_5_NUM174 (.ZN (N727), .A1 (XNOR_1_3_NUM174_OUT), .A2 (XNOR_1_4_NUM174_OUT));
      wire XNOR_1_1_NUM175_OUT, XNOR_1_2_NUM175_OUT, XNOR_1_3_NUM175_OUT, XNOR_1_4_NUM175_OUT;
      NOR2_X1 XNOR_1_1_NUM175 (.ZN (XNOR_1_1_NUM175_OUT), .A1 (N17), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM175 (.ZN (XNOR_1_2_NUM175_OUT), .A1 (GND), .A2 (N696));
      NOR2_X1 XNOR_1_3_NUM175 (.ZN (XNOR_1_3_NUM175_OUT), .A1 (XNOR_1_1_NUM175_OUT), .A2 (XNOR_1_2_NUM175_OUT));
      NOR2_X1 XNOR_1_4_NUM175 (.ZN (XNOR_1_4_NUM175_OUT), .A1 (N17), .A2 (N696));
      NOR2_X1 XNOR_1_5_NUM175 (.ZN (N728), .A1 (XNOR_1_3_NUM175_OUT), .A2 (XNOR_1_4_NUM175_OUT));
      wire XNOR_1_1_NUM176_OUT, XNOR_1_2_NUM176_OUT, XNOR_1_3_NUM176_OUT, XNOR_1_4_NUM176_OUT;
      NOR2_X1 XNOR_1_1_NUM176 (.ZN (XNOR_1_1_NUM176_OUT), .A1 (N21), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM176 (.ZN (XNOR_1_2_NUM176_OUT), .A1 (GND), .A2 (N697));
      NOR2_X1 XNOR_1_3_NUM176 (.ZN (XNOR_1_3_NUM176_OUT), .A1 (XNOR_1_1_NUM176_OUT), .A2 (XNOR_1_2_NUM176_OUT));
      NOR2_X1 XNOR_1_4_NUM176 (.ZN (XNOR_1_4_NUM176_OUT), .A1 (N21), .A2 (N697));
      NOR2_X1 XNOR_1_5_NUM176 (.ZN (N729), .A1 (XNOR_1_3_NUM176_OUT), .A2 (XNOR_1_4_NUM176_OUT));
      wire XNOR_1_1_NUM177_OUT, XNOR_1_2_NUM177_OUT, XNOR_1_3_NUM177_OUT, XNOR_1_4_NUM177_OUT;
      NOR2_X1 XNOR_1_1_NUM177 (.ZN (XNOR_1_1_NUM177_OUT), .A1 (N25), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM177 (.ZN (XNOR_1_2_NUM177_OUT), .A1 (GND), .A2 (N698));
      NOR2_X1 XNOR_1_3_NUM177 (.ZN (XNOR_1_3_NUM177_OUT), .A1 (XNOR_1_1_NUM177_OUT), .A2 (XNOR_1_2_NUM177_OUT));
      NOR2_X1 XNOR_1_4_NUM177 (.ZN (XNOR_1_4_NUM177_OUT), .A1 (N25), .A2 (N698));
      NOR2_X1 XNOR_1_5_NUM177 (.ZN (N730), .A1 (XNOR_1_3_NUM177_OUT), .A2 (XNOR_1_4_NUM177_OUT));
      wire XNOR_1_1_NUM178_OUT, XNOR_1_2_NUM178_OUT, XNOR_1_3_NUM178_OUT, XNOR_1_4_NUM178_OUT;
      NOR2_X1 XNOR_1_1_NUM178 (.ZN (XNOR_1_1_NUM178_OUT), .A1 (N29), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM178 (.ZN (XNOR_1_2_NUM178_OUT), .A1 (GND), .A2 (N699));
      NOR2_X1 XNOR_1_3_NUM178 (.ZN (XNOR_1_3_NUM178_OUT), .A1 (XNOR_1_1_NUM178_OUT), .A2 (XNOR_1_2_NUM178_OUT));
      NOR2_X1 XNOR_1_4_NUM178 (.ZN (XNOR_1_4_NUM178_OUT), .A1 (N29), .A2 (N699));
      NOR2_X1 XNOR_1_5_NUM178 (.ZN (N731), .A1 (XNOR_1_3_NUM178_OUT), .A2 (XNOR_1_4_NUM178_OUT));
      wire XNOR_1_1_NUM179_OUT, XNOR_1_2_NUM179_OUT, XNOR_1_3_NUM179_OUT, XNOR_1_4_NUM179_OUT;
      NOR2_X1 XNOR_1_1_NUM179 (.ZN (XNOR_1_1_NUM179_OUT), .A1 (N33), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM179 (.ZN (XNOR_1_2_NUM179_OUT), .A1 (GND), .A2 (N700));
      NOR2_X1 XNOR_1_3_NUM179 (.ZN (XNOR_1_3_NUM179_OUT), .A1 (XNOR_1_1_NUM179_OUT), .A2 (XNOR_1_2_NUM179_OUT));
      NOR2_X1 XNOR_1_4_NUM179 (.ZN (XNOR_1_4_NUM179_OUT), .A1 (N33), .A2 (N700));
      NOR2_X1 XNOR_1_5_NUM179 (.ZN (N732), .A1 (XNOR_1_3_NUM179_OUT), .A2 (XNOR_1_4_NUM179_OUT));
      wire XNOR_1_1_NUM180_OUT, XNOR_1_2_NUM180_OUT, XNOR_1_3_NUM180_OUT, XNOR_1_4_NUM180_OUT;
      NOR2_X1 XNOR_1_1_NUM180 (.ZN (XNOR_1_1_NUM180_OUT), .A1 (N37), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM180 (.ZN (XNOR_1_2_NUM180_OUT), .A1 (GND), .A2 (N701));
      NOR2_X1 XNOR_1_3_NUM180 (.ZN (XNOR_1_3_NUM180_OUT), .A1 (XNOR_1_1_NUM180_OUT), .A2 (XNOR_1_2_NUM180_OUT));
      NOR2_X1 XNOR_1_4_NUM180 (.ZN (XNOR_1_4_NUM180_OUT), .A1 (N37), .A2 (N701));
      NOR2_X1 XNOR_1_5_NUM180 (.ZN (N733), .A1 (XNOR_1_3_NUM180_OUT), .A2 (XNOR_1_4_NUM180_OUT));
      wire XNOR_1_1_NUM181_OUT, XNOR_1_2_NUM181_OUT, XNOR_1_3_NUM181_OUT, XNOR_1_4_NUM181_OUT;
      NOR2_X1 XNOR_1_1_NUM181 (.ZN (XNOR_1_1_NUM181_OUT), .A1 (N41), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM181 (.ZN (XNOR_1_2_NUM181_OUT), .A1 (GND), .A2 (N702));
      NOR2_X1 XNOR_1_3_NUM181 (.ZN (XNOR_1_3_NUM181_OUT), .A1 (XNOR_1_1_NUM181_OUT), .A2 (XNOR_1_2_NUM181_OUT));
      NOR2_X1 XNOR_1_4_NUM181 (.ZN (XNOR_1_4_NUM181_OUT), .A1 (N41), .A2 (N702));
      NOR2_X1 XNOR_1_5_NUM181 (.ZN (N734), .A1 (XNOR_1_3_NUM181_OUT), .A2 (XNOR_1_4_NUM181_OUT));
      wire XNOR_1_1_NUM182_OUT, XNOR_1_2_NUM182_OUT, XNOR_1_3_NUM182_OUT, XNOR_1_4_NUM182_OUT;
      NOR2_X1 XNOR_1_1_NUM182 (.ZN (XNOR_1_1_NUM182_OUT), .A1 (N45), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM182 (.ZN (XNOR_1_2_NUM182_OUT), .A1 (GND), .A2 (N703));
      NOR2_X1 XNOR_1_3_NUM182 (.ZN (XNOR_1_3_NUM182_OUT), .A1 (XNOR_1_1_NUM182_OUT), .A2 (XNOR_1_2_NUM182_OUT));
      NOR2_X1 XNOR_1_4_NUM182 (.ZN (XNOR_1_4_NUM182_OUT), .A1 (N45), .A2 (N703));
      NOR2_X1 XNOR_1_5_NUM182 (.ZN (N735), .A1 (XNOR_1_3_NUM182_OUT), .A2 (XNOR_1_4_NUM182_OUT));
      wire XNOR_1_1_NUM183_OUT, XNOR_1_2_NUM183_OUT, XNOR_1_3_NUM183_OUT, XNOR_1_4_NUM183_OUT;
      NOR2_X1 XNOR_1_1_NUM183 (.ZN (XNOR_1_1_NUM183_OUT), .A1 (N49), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM183 (.ZN (XNOR_1_2_NUM183_OUT), .A1 (GND), .A2 (N704));
      NOR2_X1 XNOR_1_3_NUM183 (.ZN (XNOR_1_3_NUM183_OUT), .A1 (XNOR_1_1_NUM183_OUT), .A2 (XNOR_1_2_NUM183_OUT));
      NOR2_X1 XNOR_1_4_NUM183 (.ZN (XNOR_1_4_NUM183_OUT), .A1 (N49), .A2 (N704));
      NOR2_X1 XNOR_1_5_NUM183 (.ZN (N736), .A1 (XNOR_1_3_NUM183_OUT), .A2 (XNOR_1_4_NUM183_OUT));
      wire XNOR_1_1_NUM184_OUT, XNOR_1_2_NUM184_OUT, XNOR_1_3_NUM184_OUT, XNOR_1_4_NUM184_OUT;
      NOR2_X1 XNOR_1_1_NUM184 (.ZN (XNOR_1_1_NUM184_OUT), .A1 (N53), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM184 (.ZN (XNOR_1_2_NUM184_OUT), .A1 (GND), .A2 (N705));
      NOR2_X1 XNOR_1_3_NUM184 (.ZN (XNOR_1_3_NUM184_OUT), .A1 (XNOR_1_1_NUM184_OUT), .A2 (XNOR_1_2_NUM184_OUT));
      NOR2_X1 XNOR_1_4_NUM184 (.ZN (XNOR_1_4_NUM184_OUT), .A1 (N53), .A2 (N705));
      NOR2_X1 XNOR_1_5_NUM184 (.ZN (N737), .A1 (XNOR_1_3_NUM184_OUT), .A2 (XNOR_1_4_NUM184_OUT));
      wire XNOR_1_1_NUM185_OUT, XNOR_1_2_NUM185_OUT, XNOR_1_3_NUM185_OUT, XNOR_1_4_NUM185_OUT;
      NOR2_X1 XNOR_1_1_NUM185 (.ZN (XNOR_1_1_NUM185_OUT), .A1 (N57), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM185 (.ZN (XNOR_1_2_NUM185_OUT), .A1 (GND), .A2 (N706));
      NOR2_X1 XNOR_1_3_NUM185 (.ZN (XNOR_1_3_NUM185_OUT), .A1 (XNOR_1_1_NUM185_OUT), .A2 (XNOR_1_2_NUM185_OUT));
      NOR2_X1 XNOR_1_4_NUM185 (.ZN (XNOR_1_4_NUM185_OUT), .A1 (N57), .A2 (N706));
      NOR2_X1 XNOR_1_5_NUM185 (.ZN (N738), .A1 (XNOR_1_3_NUM185_OUT), .A2 (XNOR_1_4_NUM185_OUT));
      wire XNOR_1_1_NUM186_OUT, XNOR_1_2_NUM186_OUT, XNOR_1_3_NUM186_OUT, XNOR_1_4_NUM186_OUT;
      NOR2_X1 XNOR_1_1_NUM186 (.ZN (XNOR_1_1_NUM186_OUT), .A1 (N61), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM186 (.ZN (XNOR_1_2_NUM186_OUT), .A1 (GND), .A2 (N707));
      NOR2_X1 XNOR_1_3_NUM186 (.ZN (XNOR_1_3_NUM186_OUT), .A1 (XNOR_1_1_NUM186_OUT), .A2 (XNOR_1_2_NUM186_OUT));
      NOR2_X1 XNOR_1_4_NUM186 (.ZN (XNOR_1_4_NUM186_OUT), .A1 (N61), .A2 (N707));
      NOR2_X1 XNOR_1_5_NUM186 (.ZN (N739), .A1 (XNOR_1_3_NUM186_OUT), .A2 (XNOR_1_4_NUM186_OUT));
      wire XNOR_1_1_NUM187_OUT, XNOR_1_2_NUM187_OUT, XNOR_1_3_NUM187_OUT, XNOR_1_4_NUM187_OUT;
      NOR2_X1 XNOR_1_1_NUM187 (.ZN (XNOR_1_1_NUM187_OUT), .A1 (N65), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM187 (.ZN (XNOR_1_2_NUM187_OUT), .A1 (GND), .A2 (N708));
      NOR2_X1 XNOR_1_3_NUM187 (.ZN (XNOR_1_3_NUM187_OUT), .A1 (XNOR_1_1_NUM187_OUT), .A2 (XNOR_1_2_NUM187_OUT));
      NOR2_X1 XNOR_1_4_NUM187 (.ZN (XNOR_1_4_NUM187_OUT), .A1 (N65), .A2 (N708));
      NOR2_X1 XNOR_1_5_NUM187 (.ZN (N740), .A1 (XNOR_1_3_NUM187_OUT), .A2 (XNOR_1_4_NUM187_OUT));
      wire XNOR_1_1_NUM188_OUT, XNOR_1_2_NUM188_OUT, XNOR_1_3_NUM188_OUT, XNOR_1_4_NUM188_OUT;
      NOR2_X1 XNOR_1_1_NUM188 (.ZN (XNOR_1_1_NUM188_OUT), .A1 (N69), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM188 (.ZN (XNOR_1_2_NUM188_OUT), .A1 (GND), .A2 (N709));
      NOR2_X1 XNOR_1_3_NUM188 (.ZN (XNOR_1_3_NUM188_OUT), .A1 (XNOR_1_1_NUM188_OUT), .A2 (XNOR_1_2_NUM188_OUT));
      NOR2_X1 XNOR_1_4_NUM188 (.ZN (XNOR_1_4_NUM188_OUT), .A1 (N69), .A2 (N709));
      NOR2_X1 XNOR_1_5_NUM188 (.ZN (N741), .A1 (XNOR_1_3_NUM188_OUT), .A2 (XNOR_1_4_NUM188_OUT));
      wire XNOR_1_1_NUM189_OUT, XNOR_1_2_NUM189_OUT, XNOR_1_3_NUM189_OUT, XNOR_1_4_NUM189_OUT;
      NOR2_X1 XNOR_1_1_NUM189 (.ZN (XNOR_1_1_NUM189_OUT), .A1 (N73), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM189 (.ZN (XNOR_1_2_NUM189_OUT), .A1 (GND), .A2 (N710));
      NOR2_X1 XNOR_1_3_NUM189 (.ZN (XNOR_1_3_NUM189_OUT), .A1 (XNOR_1_1_NUM189_OUT), .A2 (XNOR_1_2_NUM189_OUT));
      NOR2_X1 XNOR_1_4_NUM189 (.ZN (XNOR_1_4_NUM189_OUT), .A1 (N73), .A2 (N710));
      NOR2_X1 XNOR_1_5_NUM189 (.ZN (N742), .A1 (XNOR_1_3_NUM189_OUT), .A2 (XNOR_1_4_NUM189_OUT));
      wire XNOR_1_1_NUM190_OUT, XNOR_1_2_NUM190_OUT, XNOR_1_3_NUM190_OUT, XNOR_1_4_NUM190_OUT;
      NOR2_X1 XNOR_1_1_NUM190 (.ZN (XNOR_1_1_NUM190_OUT), .A1 (N77), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM190 (.ZN (XNOR_1_2_NUM190_OUT), .A1 (GND), .A2 (N711));
      NOR2_X1 XNOR_1_3_NUM190 (.ZN (XNOR_1_3_NUM190_OUT), .A1 (XNOR_1_1_NUM190_OUT), .A2 (XNOR_1_2_NUM190_OUT));
      NOR2_X1 XNOR_1_4_NUM190 (.ZN (XNOR_1_4_NUM190_OUT), .A1 (N77), .A2 (N711));
      NOR2_X1 XNOR_1_5_NUM190 (.ZN (N743), .A1 (XNOR_1_3_NUM190_OUT), .A2 (XNOR_1_4_NUM190_OUT));
      wire XNOR_1_1_NUM191_OUT, XNOR_1_2_NUM191_OUT, XNOR_1_3_NUM191_OUT, XNOR_1_4_NUM191_OUT;
      NOR2_X1 XNOR_1_1_NUM191 (.ZN (XNOR_1_1_NUM191_OUT), .A1 (N81), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM191 (.ZN (XNOR_1_2_NUM191_OUT), .A1 (GND), .A2 (N712));
      NOR2_X1 XNOR_1_3_NUM191 (.ZN (XNOR_1_3_NUM191_OUT), .A1 (XNOR_1_1_NUM191_OUT), .A2 (XNOR_1_2_NUM191_OUT));
      NOR2_X1 XNOR_1_4_NUM191 (.ZN (XNOR_1_4_NUM191_OUT), .A1 (N81), .A2 (N712));
      NOR2_X1 XNOR_1_5_NUM191 (.ZN (N744), .A1 (XNOR_1_3_NUM191_OUT), .A2 (XNOR_1_4_NUM191_OUT));
      wire XNOR_1_1_NUM192_OUT, XNOR_1_2_NUM192_OUT, XNOR_1_3_NUM192_OUT, XNOR_1_4_NUM192_OUT;
      NOR2_X1 XNOR_1_1_NUM192 (.ZN (XNOR_1_1_NUM192_OUT), .A1 (N85), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM192 (.ZN (XNOR_1_2_NUM192_OUT), .A1 (GND), .A2 (N713));
      NOR2_X1 XNOR_1_3_NUM192 (.ZN (XNOR_1_3_NUM192_OUT), .A1 (XNOR_1_1_NUM192_OUT), .A2 (XNOR_1_2_NUM192_OUT));
      NOR2_X1 XNOR_1_4_NUM192 (.ZN (XNOR_1_4_NUM192_OUT), .A1 (N85), .A2 (N713));
      NOR2_X1 XNOR_1_5_NUM192 (.ZN (N745), .A1 (XNOR_1_3_NUM192_OUT), .A2 (XNOR_1_4_NUM192_OUT));
      wire XNOR_1_1_NUM193_OUT, XNOR_1_2_NUM193_OUT, XNOR_1_3_NUM193_OUT, XNOR_1_4_NUM193_OUT;
      NOR2_X1 XNOR_1_1_NUM193 (.ZN (XNOR_1_1_NUM193_OUT), .A1 (N89), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM193 (.ZN (XNOR_1_2_NUM193_OUT), .A1 (GND), .A2 (N714));
      NOR2_X1 XNOR_1_3_NUM193 (.ZN (XNOR_1_3_NUM193_OUT), .A1 (XNOR_1_1_NUM193_OUT), .A2 (XNOR_1_2_NUM193_OUT));
      NOR2_X1 XNOR_1_4_NUM193 (.ZN (XNOR_1_4_NUM193_OUT), .A1 (N89), .A2 (N714));
      NOR2_X1 XNOR_1_5_NUM193 (.ZN (N746), .A1 (XNOR_1_3_NUM193_OUT), .A2 (XNOR_1_4_NUM193_OUT));
      wire XNOR_1_1_NUM194_OUT, XNOR_1_2_NUM194_OUT, XNOR_1_3_NUM194_OUT, XNOR_1_4_NUM194_OUT;
      NOR2_X1 XNOR_1_1_NUM194 (.ZN (XNOR_1_1_NUM194_OUT), .A1 (N93), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM194 (.ZN (XNOR_1_2_NUM194_OUT), .A1 (GND), .A2 (N715));
      NOR2_X1 XNOR_1_3_NUM194 (.ZN (XNOR_1_3_NUM194_OUT), .A1 (XNOR_1_1_NUM194_OUT), .A2 (XNOR_1_2_NUM194_OUT));
      NOR2_X1 XNOR_1_4_NUM194 (.ZN (XNOR_1_4_NUM194_OUT), .A1 (N93), .A2 (N715));
      NOR2_X1 XNOR_1_5_NUM194 (.ZN (N747), .A1 (XNOR_1_3_NUM194_OUT), .A2 (XNOR_1_4_NUM194_OUT));
      wire XNOR_1_1_NUM195_OUT, XNOR_1_2_NUM195_OUT, XNOR_1_3_NUM195_OUT, XNOR_1_4_NUM195_OUT;
      NOR2_X1 XNOR_1_1_NUM195 (.ZN (XNOR_1_1_NUM195_OUT), .A1 (N97), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM195 (.ZN (XNOR_1_2_NUM195_OUT), .A1 (GND), .A2 (N716));
      NOR2_X1 XNOR_1_3_NUM195 (.ZN (XNOR_1_3_NUM195_OUT), .A1 (XNOR_1_1_NUM195_OUT), .A2 (XNOR_1_2_NUM195_OUT));
      NOR2_X1 XNOR_1_4_NUM195 (.ZN (XNOR_1_4_NUM195_OUT), .A1 (N97), .A2 (N716));
      NOR2_X1 XNOR_1_5_NUM195 (.ZN (N748), .A1 (XNOR_1_3_NUM195_OUT), .A2 (XNOR_1_4_NUM195_OUT));
      wire XNOR_1_1_NUM196_OUT, XNOR_1_2_NUM196_OUT, XNOR_1_3_NUM196_OUT, XNOR_1_4_NUM196_OUT;
      NOR2_X1 XNOR_1_1_NUM196 (.ZN (XNOR_1_1_NUM196_OUT), .A1 (N101), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM196 (.ZN (XNOR_1_2_NUM196_OUT), .A1 (GND), .A2 (N717));
      NOR2_X1 XNOR_1_3_NUM196 (.ZN (XNOR_1_3_NUM196_OUT), .A1 (XNOR_1_1_NUM196_OUT), .A2 (XNOR_1_2_NUM196_OUT));
      NOR2_X1 XNOR_1_4_NUM196 (.ZN (XNOR_1_4_NUM196_OUT), .A1 (N101), .A2 (N717));
      NOR2_X1 XNOR_1_5_NUM196 (.ZN (N749), .A1 (XNOR_1_3_NUM196_OUT), .A2 (XNOR_1_4_NUM196_OUT));
      wire XNOR_1_1_NUM197_OUT, XNOR_1_2_NUM197_OUT, XNOR_1_3_NUM197_OUT, XNOR_1_4_NUM197_OUT;
      NOR2_X1 XNOR_1_1_NUM197 (.ZN (XNOR_1_1_NUM197_OUT), .A1 (N105), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM197 (.ZN (XNOR_1_2_NUM197_OUT), .A1 (GND), .A2 (N718));
      NOR2_X1 XNOR_1_3_NUM197 (.ZN (XNOR_1_3_NUM197_OUT), .A1 (XNOR_1_1_NUM197_OUT), .A2 (XNOR_1_2_NUM197_OUT));
      NOR2_X1 XNOR_1_4_NUM197 (.ZN (XNOR_1_4_NUM197_OUT), .A1 (N105), .A2 (N718));
      NOR2_X1 XNOR_1_5_NUM197 (.ZN (N750), .A1 (XNOR_1_3_NUM197_OUT), .A2 (XNOR_1_4_NUM197_OUT));
      wire XNOR_1_1_NUM198_OUT, XNOR_1_2_NUM198_OUT, XNOR_1_3_NUM198_OUT, XNOR_1_4_NUM198_OUT;
      NOR2_X1 XNOR_1_1_NUM198 (.ZN (XNOR_1_1_NUM198_OUT), .A1 (N109), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM198 (.ZN (XNOR_1_2_NUM198_OUT), .A1 (GND), .A2 (N719));
      NOR2_X1 XNOR_1_3_NUM198 (.ZN (XNOR_1_3_NUM198_OUT), .A1 (XNOR_1_1_NUM198_OUT), .A2 (XNOR_1_2_NUM198_OUT));
      NOR2_X1 XNOR_1_4_NUM198 (.ZN (XNOR_1_4_NUM198_OUT), .A1 (N109), .A2 (N719));
      NOR2_X1 XNOR_1_5_NUM198 (.ZN (N751), .A1 (XNOR_1_3_NUM198_OUT), .A2 (XNOR_1_4_NUM198_OUT));
      wire XNOR_1_1_NUM199_OUT, XNOR_1_2_NUM199_OUT, XNOR_1_3_NUM199_OUT, XNOR_1_4_NUM199_OUT;
      NOR2_X1 XNOR_1_1_NUM199 (.ZN (XNOR_1_1_NUM199_OUT), .A1 (N113), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM199 (.ZN (XNOR_1_2_NUM199_OUT), .A1 (GND), .A2 (N720));
      NOR2_X1 XNOR_1_3_NUM199 (.ZN (XNOR_1_3_NUM199_OUT), .A1 (XNOR_1_1_NUM199_OUT), .A2 (XNOR_1_2_NUM199_OUT));
      NOR2_X1 XNOR_1_4_NUM199 (.ZN (XNOR_1_4_NUM199_OUT), .A1 (N113), .A2 (N720));
      NOR2_X1 XNOR_1_5_NUM199 (.ZN (N752), .A1 (XNOR_1_3_NUM199_OUT), .A2 (XNOR_1_4_NUM199_OUT));
      wire XNOR_1_1_NUM200_OUT, XNOR_1_2_NUM200_OUT, XNOR_1_3_NUM200_OUT, XNOR_1_4_NUM200_OUT;
      NOR2_X1 XNOR_1_1_NUM200 (.ZN (XNOR_1_1_NUM200_OUT), .A1 (N117), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM200 (.ZN (XNOR_1_2_NUM200_OUT), .A1 (GND), .A2 (N721));
      NOR2_X1 XNOR_1_3_NUM200 (.ZN (XNOR_1_3_NUM200_OUT), .A1 (XNOR_1_1_NUM200_OUT), .A2 (XNOR_1_2_NUM200_OUT));
      NOR2_X1 XNOR_1_4_NUM200 (.ZN (XNOR_1_4_NUM200_OUT), .A1 (N117), .A2 (N721));
      NOR2_X1 XNOR_1_5_NUM200 (.ZN (N753), .A1 (XNOR_1_3_NUM200_OUT), .A2 (XNOR_1_4_NUM200_OUT));
      wire XNOR_1_1_NUM201_OUT, XNOR_1_2_NUM201_OUT, XNOR_1_3_NUM201_OUT, XNOR_1_4_NUM201_OUT;
      NOR2_X1 XNOR_1_1_NUM201 (.ZN (XNOR_1_1_NUM201_OUT), .A1 (N121), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM201 (.ZN (XNOR_1_2_NUM201_OUT), .A1 (GND), .A2 (N722));
      NOR2_X1 XNOR_1_3_NUM201 (.ZN (XNOR_1_3_NUM201_OUT), .A1 (XNOR_1_1_NUM201_OUT), .A2 (XNOR_1_2_NUM201_OUT));
      NOR2_X1 XNOR_1_4_NUM201 (.ZN (XNOR_1_4_NUM201_OUT), .A1 (N121), .A2 (N722));
      NOR2_X1 XNOR_1_5_NUM201 (.ZN (N754), .A1 (XNOR_1_3_NUM201_OUT), .A2 (XNOR_1_4_NUM201_OUT));
      wire XNOR_1_1_NUM202_OUT, XNOR_1_2_NUM202_OUT, XNOR_1_3_NUM202_OUT, XNOR_1_4_NUM202_OUT;
      NOR2_X1 XNOR_1_1_NUM202 (.ZN (XNOR_1_1_NUM202_OUT), .A1 (N125), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM202 (.ZN (XNOR_1_2_NUM202_OUT), .A1 (GND), .A2 (N723));
      NOR2_X1 XNOR_1_3_NUM202 (.ZN (XNOR_1_3_NUM202_OUT), .A1 (XNOR_1_1_NUM202_OUT), .A2 (XNOR_1_2_NUM202_OUT));
      NOR2_X1 XNOR_1_4_NUM202 (.ZN (XNOR_1_4_NUM202_OUT), .A1 (N125), .A2 (N723));
      NOR2_X1 XNOR_1_5_NUM202 (.ZN (N755), .A1 (XNOR_1_3_NUM202_OUT), .A2 (XNOR_1_4_NUM202_OUT));


      wire XNOR_1_1_N724_TERMINATION_OUT, XNOR_1_2_N724_TERMINATION_OUT;
      NOR2_X1 XNOR_1_1_N724_TERMINATION (.ZN (XNOR_1_1_N724_TERMINATION_OUT), .A1 (N724), .A2 (GND));
      NOR2_X1 XNOR_1_2_N724_TERMINATION (.ZN (N724_TERMINATION), .A1 (XNOR_1_1_N724_TERMINATION_OUT), .A2 (XNOR_1_2_N724_TERMINATION_OUT));

      wire XNOR_1_1_N725_TERMINATION_OUT, XNOR_1_2_N725_TERMINATION_OUT;
      NOR2_X1 XNOR_1_1_N725_TERMINATION (.ZN (XNOR_1_1_N725_TERMINATION_OUT), .A1 (N725), .A2 (GND));
      NOR2_X1 XNOR_1_2_N725_TERMINATION (.ZN (N725_TERMINATION), .A1 (XNOR_1_1_N725_TERMINATION_OUT), .A2 (XNOR_1_2_N725_TERMINATION_OUT));

      wire XNOR_1_1_N726_TERMINATION_OUT, XNOR_1_2_N726_TERMINATION_OUT;
      NOR2_X1 XNOR_1_1_N726_TERMINATION (.ZN (XNOR_1_1_N726_TERMINATION_OUT), .A1 (N726), .A2 (GND));
      NOR2_X1 XNOR_1_2_N726_TERMINATION (.ZN (N726_TERMINATION), .A1 (XNOR_1_1_N726_TERMINATION_OUT), .A2 (XNOR_1_2_N726_TERMINATION_OUT));

      wire XNOR_1_1_N727_TERMINATION_OUT, XNOR_1_2_N727_TERMINATION_OUT;
      NOR2_X1 XNOR_1_1_N727_TERMINATION (.ZN (XNOR_1_1_N727_TERMINATION_OUT), .A1 (N727), .A2 (GND));
      NOR2_X1 XNOR_1_2_N727_TERMINATION (.ZN (N727_TERMINATION), .A1 (XNOR_1_1_N727_TERMINATION_OUT), .A2 (XNOR_1_2_N727_TERMINATION_OUT));

      wire XNOR_1_1_N728_TERMINATION_OUT, XNOR_1_2_N728_TERMINATION_OUT;
      NOR2_X1 XNOR_1_1_N728_TERMINATION (.ZN (XNOR_1_1_N728_TERMINATION_OUT), .A1 (N728), .A2 (GND));
      NOR2_X1 XNOR_1_2_N728_TERMINATION (.ZN (N728_TERMINATION), .A1 (XNOR_1_1_N728_TERMINATION_OUT), .A2 (XNOR_1_2_N728_TERMINATION_OUT));

      wire XNOR_1_1_N729_TERMINATION_OUT, XNOR_1_2_N729_TERMINATION_OUT;
      NOR2_X1 XNOR_1_1_N729_TERMINATION (.ZN (XNOR_1_1_N729_TERMINATION_OUT), .A1 (N729), .A2 (GND));
      NOR2_X1 XNOR_1_2_N729_TERMINATION (.ZN (N729_TERMINATION), .A1 (XNOR_1_1_N729_TERMINATION_OUT), .A2 (XNOR_1_2_N729_TERMINATION_OUT));

      wire XNOR_1_1_N730_TERMINATION_OUT, XNOR_1_2_N730_TERMINATION_OUT;
      NOR2_X1 XNOR_1_1_N730_TERMINATION (.ZN (XNOR_1_1_N730_TERMINATION_OUT), .A1 (N730), .A2 (GND));
      NOR2_X1 XNOR_1_2_N730_TERMINATION (.ZN (N730_TERMINATION), .A1 (XNOR_1_1_N730_TERMINATION_OUT), .A2 (XNOR_1_2_N730_TERMINATION_OUT));

      wire XNOR_1_1_N731_TERMINATION_OUT, XNOR_1_2_N731_TERMINATION_OUT;
      NOR2_X1 XNOR_1_1_N731_TERMINATION (.ZN (XNOR_1_1_N731_TERMINATION_OUT), .A1 (N731), .A2 (GND));
      NOR2_X1 XNOR_1_2_N731_TERMINATION (.ZN (N731_TERMINATION), .A1 (XNOR_1_1_N731_TERMINATION_OUT), .A2 (XNOR_1_2_N731_TERMINATION_OUT));

      wire XNOR_1_1_N732_TERMINATION_OUT, XNOR_1_2_N732_TERMINATION_OUT;
      NOR2_X1 XNOR_1_1_N732_TERMINATION (.ZN (XNOR_1_1_N732_TERMINATION_OUT), .A1 (N732), .A2 (GND));
      NOR2_X1 XNOR_1_2_N732_TERMINATION (.ZN (N732_TERMINATION), .A1 (XNOR_1_1_N732_TERMINATION_OUT), .A2 (XNOR_1_2_N732_TERMINATION_OUT));

      wire XNOR_1_1_N733_TERMINATION_OUT, XNOR_1_2_N733_TERMINATION_OUT;
      NOR2_X1 XNOR_1_1_N733_TERMINATION (.ZN (XNOR_1_1_N733_TERMINATION_OUT), .A1 (N733), .A2 (GND));
      NOR2_X1 XNOR_1_2_N733_TERMINATION (.ZN (N733_TERMINATION), .A1 (XNOR_1_1_N733_TERMINATION_OUT), .A2 (XNOR_1_2_N733_TERMINATION_OUT));

      wire XNOR_1_1_N734_TERMINATION_OUT, XNOR_1_2_N734_TERMINATION_OUT;
      NOR2_X1 XNOR_1_1_N734_TERMINATION (.ZN (XNOR_1_1_N734_TERMINATION_OUT), .A1 (N734), .A2 (GND));
      NOR2_X1 XNOR_1_2_N734_TERMINATION (.ZN (N734_TERMINATION), .A1 (XNOR_1_1_N734_TERMINATION_OUT), .A2 (XNOR_1_2_N734_TERMINATION_OUT));

      wire XNOR_1_1_N735_TERMINATION_OUT, XNOR_1_2_N735_TERMINATION_OUT;
      NOR2_X1 XNOR_1_1_N735_TERMINATION (.ZN (XNOR_1_1_N735_TERMINATION_OUT), .A1 (N735), .A2 (GND));
      NOR2_X1 XNOR_1_2_N735_TERMINATION (.ZN (N735_TERMINATION), .A1 (XNOR_1_1_N735_TERMINATION_OUT), .A2 (XNOR_1_2_N735_TERMINATION_OUT));

      wire XNOR_1_1_N736_TERMINATION_OUT, XNOR_1_2_N736_TERMINATION_OUT;
      NOR2_X1 XNOR_1_1_N736_TERMINATION (.ZN (XNOR_1_1_N736_TERMINATION_OUT), .A1 (N736), .A2 (GND));
      NOR2_X1 XNOR_1_2_N736_TERMINATION (.ZN (N736_TERMINATION), .A1 (XNOR_1_1_N736_TERMINATION_OUT), .A2 (XNOR_1_2_N736_TERMINATION_OUT));

      wire XNOR_1_1_N737_TERMINATION_OUT, XNOR_1_2_N737_TERMINATION_OUT;
      NOR2_X1 XNOR_1_1_N737_TERMINATION (.ZN (XNOR_1_1_N737_TERMINATION_OUT), .A1 (N737), .A2 (GND));
      NOR2_X1 XNOR_1_2_N737_TERMINATION (.ZN (N737_TERMINATION), .A1 (XNOR_1_1_N737_TERMINATION_OUT), .A2 (XNOR_1_2_N737_TERMINATION_OUT));

      wire XNOR_1_1_N738_TERMINATION_OUT, XNOR_1_2_N738_TERMINATION_OUT;
      NOR2_X1 XNOR_1_1_N738_TERMINATION (.ZN (XNOR_1_1_N738_TERMINATION_OUT), .A1 (N738), .A2 (GND));
      NOR2_X1 XNOR_1_2_N738_TERMINATION (.ZN (N738_TERMINATION), .A1 (XNOR_1_1_N738_TERMINATION_OUT), .A2 (XNOR_1_2_N738_TERMINATION_OUT));

      wire XNOR_1_1_N739_TERMINATION_OUT, XNOR_1_2_N739_TERMINATION_OUT;
      NOR2_X1 XNOR_1_1_N739_TERMINATION (.ZN (XNOR_1_1_N739_TERMINATION_OUT), .A1 (N739), .A2 (GND));
      NOR2_X1 XNOR_1_2_N739_TERMINATION (.ZN (N739_TERMINATION), .A1 (XNOR_1_1_N739_TERMINATION_OUT), .A2 (XNOR_1_2_N739_TERMINATION_OUT));

      wire XNOR_1_1_N740_TERMINATION_OUT, XNOR_1_2_N740_TERMINATION_OUT;
      NOR2_X1 XNOR_1_1_N740_TERMINATION (.ZN (XNOR_1_1_N740_TERMINATION_OUT), .A1 (N740), .A2 (GND));
      NOR2_X1 XNOR_1_2_N740_TERMINATION (.ZN (N740_TERMINATION), .A1 (XNOR_1_1_N740_TERMINATION_OUT), .A2 (XNOR_1_2_N740_TERMINATION_OUT));

      wire XNOR_1_1_N741_TERMINATION_OUT, XNOR_1_2_N741_TERMINATION_OUT;
      NOR2_X1 XNOR_1_1_N741_TERMINATION (.ZN (XNOR_1_1_N741_TERMINATION_OUT), .A1 (N741), .A2 (GND));
      NOR2_X1 XNOR_1_2_N741_TERMINATION (.ZN (N741_TERMINATION), .A1 (XNOR_1_1_N741_TERMINATION_OUT), .A2 (XNOR_1_2_N741_TERMINATION_OUT));

      wire XNOR_1_1_N742_TERMINATION_OUT, XNOR_1_2_N742_TERMINATION_OUT;
      NOR2_X1 XNOR_1_1_N742_TERMINATION (.ZN (XNOR_1_1_N742_TERMINATION_OUT), .A1 (N742), .A2 (GND));
      NOR2_X1 XNOR_1_2_N742_TERMINATION (.ZN (N742_TERMINATION), .A1 (XNOR_1_1_N742_TERMINATION_OUT), .A2 (XNOR_1_2_N742_TERMINATION_OUT));

      wire XNOR_1_1_N743_TERMINATION_OUT, XNOR_1_2_N743_TERMINATION_OUT;
      NOR2_X1 XNOR_1_1_N743_TERMINATION (.ZN (XNOR_1_1_N743_TERMINATION_OUT), .A1 (N743), .A2 (GND));
      NOR2_X1 XNOR_1_2_N743_TERMINATION (.ZN (N743_TERMINATION), .A1 (XNOR_1_1_N743_TERMINATION_OUT), .A2 (XNOR_1_2_N743_TERMINATION_OUT));

      wire XNOR_1_1_N744_TERMINATION_OUT, XNOR_1_2_N744_TERMINATION_OUT;
      NOR2_X1 XNOR_1_1_N744_TERMINATION (.ZN (XNOR_1_1_N744_TERMINATION_OUT), .A1 (N744), .A2 (GND));
      NOR2_X1 XNOR_1_2_N744_TERMINATION (.ZN (N744_TERMINATION), .A1 (XNOR_1_1_N744_TERMINATION_OUT), .A2 (XNOR_1_2_N744_TERMINATION_OUT));

      wire XNOR_1_1_N745_TERMINATION_OUT, XNOR_1_2_N745_TERMINATION_OUT;
      NOR2_X1 XNOR_1_1_N745_TERMINATION (.ZN (XNOR_1_1_N745_TERMINATION_OUT), .A1 (N745), .A2 (GND));
      NOR2_X1 XNOR_1_2_N745_TERMINATION (.ZN (N745_TERMINATION), .A1 (XNOR_1_1_N745_TERMINATION_OUT), .A2 (XNOR_1_2_N745_TERMINATION_OUT));

      wire XNOR_1_1_N746_TERMINATION_OUT, XNOR_1_2_N746_TERMINATION_OUT;
      NOR2_X1 XNOR_1_1_N746_TERMINATION (.ZN (XNOR_1_1_N746_TERMINATION_OUT), .A1 (N746), .A2 (GND));
      NOR2_X1 XNOR_1_2_N746_TERMINATION (.ZN (N746_TERMINATION), .A1 (XNOR_1_1_N746_TERMINATION_OUT), .A2 (XNOR_1_2_N746_TERMINATION_OUT));

      wire XNOR_1_1_N747_TERMINATION_OUT, XNOR_1_2_N747_TERMINATION_OUT;
      NOR2_X1 XNOR_1_1_N747_TERMINATION (.ZN (XNOR_1_1_N747_TERMINATION_OUT), .A1 (N747), .A2 (GND));
      NOR2_X1 XNOR_1_2_N747_TERMINATION (.ZN (N747_TERMINATION), .A1 (XNOR_1_1_N747_TERMINATION_OUT), .A2 (XNOR_1_2_N747_TERMINATION_OUT));

      wire XNOR_1_1_N748_TERMINATION_OUT, XNOR_1_2_N748_TERMINATION_OUT;
      NOR2_X1 XNOR_1_1_N748_TERMINATION (.ZN (XNOR_1_1_N748_TERMINATION_OUT), .A1 (N748), .A2 (GND));
      NOR2_X1 XNOR_1_2_N748_TERMINATION (.ZN (N748_TERMINATION), .A1 (XNOR_1_1_N748_TERMINATION_OUT), .A2 (XNOR_1_2_N748_TERMINATION_OUT));

      wire XNOR_1_1_N749_TERMINATION_OUT, XNOR_1_2_N749_TERMINATION_OUT;
      NOR2_X1 XNOR_1_1_N749_TERMINATION (.ZN (XNOR_1_1_N749_TERMINATION_OUT), .A1 (N749), .A2 (GND));
      NOR2_X1 XNOR_1_2_N749_TERMINATION (.ZN (N749_TERMINATION), .A1 (XNOR_1_1_N749_TERMINATION_OUT), .A2 (XNOR_1_2_N749_TERMINATION_OUT));

      wire XNOR_1_1_N750_TERMINATION_OUT, XNOR_1_2_N750_TERMINATION_OUT;
      NOR2_X1 XNOR_1_1_N750_TERMINATION (.ZN (XNOR_1_1_N750_TERMINATION_OUT), .A1 (N750), .A2 (GND));
      NOR2_X1 XNOR_1_2_N750_TERMINATION (.ZN (N750_TERMINATION), .A1 (XNOR_1_1_N750_TERMINATION_OUT), .A2 (XNOR_1_2_N750_TERMINATION_OUT));

      wire XNOR_1_1_N751_TERMINATION_OUT, XNOR_1_2_N751_TERMINATION_OUT;
      NOR2_X1 XNOR_1_1_N751_TERMINATION (.ZN (XNOR_1_1_N751_TERMINATION_OUT), .A1 (N751), .A2 (GND));
      NOR2_X1 XNOR_1_2_N751_TERMINATION (.ZN (N751_TERMINATION), .A1 (XNOR_1_1_N751_TERMINATION_OUT), .A2 (XNOR_1_2_N751_TERMINATION_OUT));

      wire XNOR_1_1_N752_TERMINATION_OUT, XNOR_1_2_N752_TERMINATION_OUT;
      NOR2_X1 XNOR_1_1_N752_TERMINATION (.ZN (XNOR_1_1_N752_TERMINATION_OUT), .A1 (N752), .A2 (GND));
      NOR2_X1 XNOR_1_2_N752_TERMINATION (.ZN (N752_TERMINATION), .A1 (XNOR_1_1_N752_TERMINATION_OUT), .A2 (XNOR_1_2_N752_TERMINATION_OUT));

      wire XNOR_1_1_N753_TERMINATION_OUT, XNOR_1_2_N753_TERMINATION_OUT;
      NOR2_X1 XNOR_1_1_N753_TERMINATION (.ZN (XNOR_1_1_N753_TERMINATION_OUT), .A1 (N753), .A2 (GND));
      NOR2_X1 XNOR_1_2_N753_TERMINATION (.ZN (N753_TERMINATION), .A1 (XNOR_1_1_N753_TERMINATION_OUT), .A2 (XNOR_1_2_N753_TERMINATION_OUT));

      wire XNOR_1_1_N754_TERMINATION_OUT, XNOR_1_2_N754_TERMINATION_OUT;
      NOR2_X1 XNOR_1_1_N754_TERMINATION (.ZN (XNOR_1_1_N754_TERMINATION_OUT), .A1 (N754), .A2 (GND));
      NOR2_X1 XNOR_1_2_N754_TERMINATION (.ZN (N754_TERMINATION), .A1 (XNOR_1_1_N754_TERMINATION_OUT), .A2 (XNOR_1_2_N754_TERMINATION_OUT));

      wire XNOR_1_1_N755_TERMINATION_OUT, XNOR_1_2_N755_TERMINATION_OUT;
      NOR2_X1 XNOR_1_1_N755_TERMINATION (.ZN (XNOR_1_1_N755_TERMINATION_OUT), .A1 (N755), .A2 (GND));
      NOR2_X1 XNOR_1_2_N755_TERMINATION (.ZN (N755_TERMINATION), .A1 (XNOR_1_1_N755_TERMINATION_OUT), .A2 (XNOR_1_2_N755_TERMINATION_OUT));


endmodule
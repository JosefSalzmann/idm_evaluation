module c432_NOR_template (N1_PWL,N4_PWL,N8_PWL,N11_PWL,N14_PWL,N17_PWL,N21_PWL,N24_PWL,N27_PWL,N30_PWL,
       N34_PWL,N37_PWL,N40_PWL,N43_PWL,N47_PWL,N50_PWL,N53_PWL,N56_PWL,N60_PWL,N63_PWL,
       N66_PWL,N69_PWL,N73_PWL,N76_PWL,N79_PWL,N82_PWL,N86_PWL,N89_PWL,N92_PWL,N95_PWL,
       N99_PWL,N102_PWL,N105_PWL,N108_PWL,N112_PWL,N115_PWL,N223_TERMINATION,N329_TERMINATION,N370_TERMINATION,N421_TERMINATION,N430_TERMINATION,N431_TERMINATION,N432_TERMINATION);

       input N1_PWL,N4_PWL,N8_PWL,N11_PWL,N14_PWL,N17_PWL,N21_PWL,N24_PWL,N27_PWL,N30_PWL,
       N34_PWL,N37_PWL,N40_PWL,N43_PWL,N47_PWL,N50_PWL,N53_PWL,N56_PWL,N60_PWL,N63_PWL,
       N66_PWL,N69_PWL,N73_PWL,N76_PWL,N79_PWL,N82_PWL,N86_PWL,N89_PWL,N92_PWL,N95_PWL,
       N99_PWL,N102_PWL,N105_PWL,N108_PWL,N112_PWL,N115_PWL;

       output N223_TERMINATION,N329_TERMINATION,N370_TERMINATION,N421_TERMINATION,N430_TERMINATION,N431_TERMINATION,N432_TERMINATION;

       wire GND = 1'b0;
       wire XNOR_1_1_N1_PULSESHAPING_OUT, XNOR_1_2_N1_PULSESHAPING_OUT, XNOR_1_3_N1_PULSESHAPING_OUT, XNOR_1_4_N1_PULSESHAPING_OUT, XNOR_1_5_N1_PULSESHAPING_OUT, XNOR_1_6_N1_PULSESHAPING_OUT;
       NOR2_X1 XNOR_1_1_N1_PULSESHAPING (.ZN (XNOR_1_1_N1_PULSESHAPING_OUT), .A1 (N1_PWL), .A2 (GND));
       NOR2_X1 XNOR_1_2_N1_PULSESHAPING (.ZN (XNOR_1_2_N1_PULSESHAPING_OUT), .A1 (XNOR_1_1_N1_PULSESHAPING_OUT), .A2 (GND));
       NOR2_X1 XNOR_1_3_N1_PULSESHAPING (.ZN (XNOR_1_3_N1_PULSESHAPING_OUT), .A1 (XNOR_1_2_N1_PULSESHAPING_OUT), .A2 (GND));
       NOR2_X1 XNOR_1_4_N1_PULSESHAPING (.ZN (XNOR_1_4_N1_PULSESHAPING_OUT), .A1 (XNOR_1_3_N1_PULSESHAPING_OUT), .A2 (GND));
       NOR2_X1 XNOR_1_5_N1_PULSESHAPING (.ZN (XNOR_1_5_N1_PULSESHAPING_OUT), .A1 (XNOR_1_4_N1_PULSESHAPING_OUT), .A2 (GND));
       NOR2_X1 XNOR_1_6_N1_PULSESHAPING (.ZN (XNOR_1_6_N1_PULSESHAPING_OUT), .A1 (XNOR_1_5_N1_PULSESHAPING_OUT), .A2 (GND));
       NOR2_X1 XNOR_1_7_N1_PULSESHAPING (.ZN (N1), .A1 (XNOR_1_6_N1_PULSESHAPING_OUT), .A2 (GND));

       wire XNOR_1_1_N4_PULSESHAPING_OUT, XNOR_1_2_N4_PULSESHAPING_OUT, XNOR_1_3_N4_PULSESHAPING_OUT, XNOR_1_4_N4_PULSESHAPING_OUT, XNOR_1_5_N4_PULSESHAPING_OUT, XNOR_1_6_N4_PULSESHAPING_OUT;
       NOR2_X1 XNOR_1_1_N4_PULSESHAPING (.ZN (XNOR_1_1_N4_PULSESHAPING_OUT), .A1 (N4_PWL), .A2 (GND));
       NOR2_X1 XNOR_1_2_N4_PULSESHAPING (.ZN (XNOR_1_2_N4_PULSESHAPING_OUT), .A1 (XNOR_1_1_N4_PULSESHAPING_OUT), .A2 (GND));
       NOR2_X1 XNOR_1_3_N4_PULSESHAPING (.ZN (XNOR_1_3_N4_PULSESHAPING_OUT), .A1 (XNOR_1_2_N4_PULSESHAPING_OUT), .A2 (GND));
       NOR2_X1 XNOR_1_4_N4_PULSESHAPING (.ZN (XNOR_1_4_N4_PULSESHAPING_OUT), .A1 (XNOR_1_3_N4_PULSESHAPING_OUT), .A2 (GND));
       NOR2_X1 XNOR_1_5_N4_PULSESHAPING (.ZN (XNOR_1_5_N4_PULSESHAPING_OUT), .A1 (XNOR_1_4_N4_PULSESHAPING_OUT), .A2 (GND));
       NOR2_X1 XNOR_1_6_N4_PULSESHAPING (.ZN (XNOR_1_6_N4_PULSESHAPING_OUT), .A1 (XNOR_1_5_N4_PULSESHAPING_OUT), .A2 (GND));
       NOR2_X1 XNOR_1_7_N4_PULSESHAPING (.ZN (N4), .A1 (XNOR_1_6_N4_PULSESHAPING_OUT), .A2 (GND));

       wire XNOR_1_1_N8_PULSESHAPING_OUT, XNOR_1_2_N8_PULSESHAPING_OUT, XNOR_1_3_N8_PULSESHAPING_OUT, XNOR_1_4_N8_PULSESHAPING_OUT, XNOR_1_5_N8_PULSESHAPING_OUT, XNOR_1_6_N8_PULSESHAPING_OUT;
       NOR2_X1 XNOR_1_1_N8_PULSESHAPING (.ZN (XNOR_1_1_N8_PULSESHAPING_OUT), .A1 (N8_PWL), .A2 (GND));
       NOR2_X1 XNOR_1_2_N8_PULSESHAPING (.ZN (XNOR_1_2_N8_PULSESHAPING_OUT), .A1 (XNOR_1_1_N8_PULSESHAPING_OUT), .A2 (GND));
       NOR2_X1 XNOR_1_3_N8_PULSESHAPING (.ZN (XNOR_1_3_N8_PULSESHAPING_OUT), .A1 (XNOR_1_2_N8_PULSESHAPING_OUT), .A2 (GND));
       NOR2_X1 XNOR_1_4_N8_PULSESHAPING (.ZN (XNOR_1_4_N8_PULSESHAPING_OUT), .A1 (XNOR_1_3_N8_PULSESHAPING_OUT), .A2 (GND));
       NOR2_X1 XNOR_1_5_N8_PULSESHAPING (.ZN (XNOR_1_5_N8_PULSESHAPING_OUT), .A1 (XNOR_1_4_N8_PULSESHAPING_OUT), .A2 (GND));
       NOR2_X1 XNOR_1_6_N8_PULSESHAPING (.ZN (XNOR_1_6_N8_PULSESHAPING_OUT), .A1 (XNOR_1_5_N8_PULSESHAPING_OUT), .A2 (GND));
       NOR2_X1 XNOR_1_7_N8_PULSESHAPING (.ZN (N8), .A1 (XNOR_1_6_N8_PULSESHAPING_OUT), .A2 (GND));

       wire XNOR_1_1_N11_PULSESHAPING_OUT, XNOR_1_2_N11_PULSESHAPING_OUT, XNOR_1_3_N11_PULSESHAPING_OUT, XNOR_1_4_N11_PULSESHAPING_OUT, XNOR_1_5_N11_PULSESHAPING_OUT, XNOR_1_6_N11_PULSESHAPING_OUT;
       NOR2_X1 XNOR_1_1_N11_PULSESHAPING (.ZN (XNOR_1_1_N11_PULSESHAPING_OUT), .A1 (N11_PWL), .A2 (GND));
       NOR2_X1 XNOR_1_2_N11_PULSESHAPING (.ZN (XNOR_1_2_N11_PULSESHAPING_OUT), .A1 (XNOR_1_1_N11_PULSESHAPING_OUT), .A2 (GND));
       NOR2_X1 XNOR_1_3_N11_PULSESHAPING (.ZN (XNOR_1_3_N11_PULSESHAPING_OUT), .A1 (XNOR_1_2_N11_PULSESHAPING_OUT), .A2 (GND));
       NOR2_X1 XNOR_1_4_N11_PULSESHAPING (.ZN (XNOR_1_4_N11_PULSESHAPING_OUT), .A1 (XNOR_1_3_N11_PULSESHAPING_OUT), .A2 (GND));
       NOR2_X1 XNOR_1_5_N11_PULSESHAPING (.ZN (XNOR_1_5_N11_PULSESHAPING_OUT), .A1 (XNOR_1_4_N11_PULSESHAPING_OUT), .A2 (GND));
       NOR2_X1 XNOR_1_6_N11_PULSESHAPING (.ZN (XNOR_1_6_N11_PULSESHAPING_OUT), .A1 (XNOR_1_5_N11_PULSESHAPING_OUT), .A2 (GND));
       NOR2_X1 XNOR_1_7_N11_PULSESHAPING (.ZN (N11), .A1 (XNOR_1_6_N11_PULSESHAPING_OUT), .A2 (GND));

       wire XNOR_1_1_N14_PULSESHAPING_OUT, XNOR_1_2_N14_PULSESHAPING_OUT, XNOR_1_3_N14_PULSESHAPING_OUT, XNOR_1_4_N14_PULSESHAPING_OUT, XNOR_1_5_N14_PULSESHAPING_OUT, XNOR_1_6_N14_PULSESHAPING_OUT;
       NOR2_X1 XNOR_1_1_N14_PULSESHAPING (.ZN (XNOR_1_1_N14_PULSESHAPING_OUT), .A1 (N14_PWL), .A2 (GND));
       NOR2_X1 XNOR_1_2_N14_PULSESHAPING (.ZN (XNOR_1_2_N14_PULSESHAPING_OUT), .A1 (XNOR_1_1_N14_PULSESHAPING_OUT), .A2 (GND));
       NOR2_X1 XNOR_1_3_N14_PULSESHAPING (.ZN (XNOR_1_3_N14_PULSESHAPING_OUT), .A1 (XNOR_1_2_N14_PULSESHAPING_OUT), .A2 (GND));
       NOR2_X1 XNOR_1_4_N14_PULSESHAPING (.ZN (XNOR_1_4_N14_PULSESHAPING_OUT), .A1 (XNOR_1_3_N14_PULSESHAPING_OUT), .A2 (GND));
       NOR2_X1 XNOR_1_5_N14_PULSESHAPING (.ZN (XNOR_1_5_N14_PULSESHAPING_OUT), .A1 (XNOR_1_4_N14_PULSESHAPING_OUT), .A2 (GND));
       NOR2_X1 XNOR_1_6_N14_PULSESHAPING (.ZN (XNOR_1_6_N14_PULSESHAPING_OUT), .A1 (XNOR_1_5_N14_PULSESHAPING_OUT), .A2 (GND));
       NOR2_X1 XNOR_1_7_N14_PULSESHAPING (.ZN (N14), .A1 (XNOR_1_6_N14_PULSESHAPING_OUT), .A2 (GND));

       wire XNOR_1_1_N17_PULSESHAPING_OUT, XNOR_1_2_N17_PULSESHAPING_OUT, XNOR_1_3_N17_PULSESHAPING_OUT, XNOR_1_4_N17_PULSESHAPING_OUT, XNOR_1_5_N17_PULSESHAPING_OUT, XNOR_1_6_N17_PULSESHAPING_OUT;
       NOR2_X1 XNOR_1_1_N17_PULSESHAPING (.ZN (XNOR_1_1_N17_PULSESHAPING_OUT), .A1 (N17_PWL), .A2 (GND));
       NOR2_X1 XNOR_1_2_N17_PULSESHAPING (.ZN (XNOR_1_2_N17_PULSESHAPING_OUT), .A1 (XNOR_1_1_N17_PULSESHAPING_OUT), .A2 (GND));
       NOR2_X1 XNOR_1_3_N17_PULSESHAPING (.ZN (XNOR_1_3_N17_PULSESHAPING_OUT), .A1 (XNOR_1_2_N17_PULSESHAPING_OUT), .A2 (GND));
       NOR2_X1 XNOR_1_4_N17_PULSESHAPING (.ZN (XNOR_1_4_N17_PULSESHAPING_OUT), .A1 (XNOR_1_3_N17_PULSESHAPING_OUT), .A2 (GND));
       NOR2_X1 XNOR_1_5_N17_PULSESHAPING (.ZN (XNOR_1_5_N17_PULSESHAPING_OUT), .A1 (XNOR_1_4_N17_PULSESHAPING_OUT), .A2 (GND));
       NOR2_X1 XNOR_1_6_N17_PULSESHAPING (.ZN (XNOR_1_6_N17_PULSESHAPING_OUT), .A1 (XNOR_1_5_N17_PULSESHAPING_OUT), .A2 (GND));
       NOR2_X1 XNOR_1_7_N17_PULSESHAPING (.ZN (N17), .A1 (XNOR_1_6_N17_PULSESHAPING_OUT), .A2 (GND));

       wire XNOR_1_1_N21_PULSESHAPING_OUT, XNOR_1_2_N21_PULSESHAPING_OUT, XNOR_1_3_N21_PULSESHAPING_OUT, XNOR_1_4_N21_PULSESHAPING_OUT, XNOR_1_5_N21_PULSESHAPING_OUT, XNOR_1_6_N21_PULSESHAPING_OUT;
       NOR2_X1 XNOR_1_1_N21_PULSESHAPING (.ZN (XNOR_1_1_N21_PULSESHAPING_OUT), .A1 (N21_PWL), .A2 (GND));
       NOR2_X1 XNOR_1_2_N21_PULSESHAPING (.ZN (XNOR_1_2_N21_PULSESHAPING_OUT), .A1 (XNOR_1_1_N21_PULSESHAPING_OUT), .A2 (GND));
       NOR2_X1 XNOR_1_3_N21_PULSESHAPING (.ZN (XNOR_1_3_N21_PULSESHAPING_OUT), .A1 (XNOR_1_2_N21_PULSESHAPING_OUT), .A2 (GND));
       NOR2_X1 XNOR_1_4_N21_PULSESHAPING (.ZN (XNOR_1_4_N21_PULSESHAPING_OUT), .A1 (XNOR_1_3_N21_PULSESHAPING_OUT), .A2 (GND));
       NOR2_X1 XNOR_1_5_N21_PULSESHAPING (.ZN (XNOR_1_5_N21_PULSESHAPING_OUT), .A1 (XNOR_1_4_N21_PULSESHAPING_OUT), .A2 (GND));
       NOR2_X1 XNOR_1_6_N21_PULSESHAPING (.ZN (XNOR_1_6_N21_PULSESHAPING_OUT), .A1 (XNOR_1_5_N21_PULSESHAPING_OUT), .A2 (GND));
       NOR2_X1 XNOR_1_7_N21_PULSESHAPING (.ZN (N21), .A1 (XNOR_1_6_N21_PULSESHAPING_OUT), .A2 (GND));

       wire XNOR_1_1_N24_PULSESHAPING_OUT, XNOR_1_2_N24_PULSESHAPING_OUT, XNOR_1_3_N24_PULSESHAPING_OUT, XNOR_1_4_N24_PULSESHAPING_OUT, XNOR_1_5_N24_PULSESHAPING_OUT, XNOR_1_6_N24_PULSESHAPING_OUT;
       NOR2_X1 XNOR_1_1_N24_PULSESHAPING (.ZN (XNOR_1_1_N24_PULSESHAPING_OUT), .A1 (N24_PWL), .A2 (GND));
       NOR2_X1 XNOR_1_2_N24_PULSESHAPING (.ZN (XNOR_1_2_N24_PULSESHAPING_OUT), .A1 (XNOR_1_1_N24_PULSESHAPING_OUT), .A2 (GND));
       NOR2_X1 XNOR_1_3_N24_PULSESHAPING (.ZN (XNOR_1_3_N24_PULSESHAPING_OUT), .A1 (XNOR_1_2_N24_PULSESHAPING_OUT), .A2 (GND));
       NOR2_X1 XNOR_1_4_N24_PULSESHAPING (.ZN (XNOR_1_4_N24_PULSESHAPING_OUT), .A1 (XNOR_1_3_N24_PULSESHAPING_OUT), .A2 (GND));
       NOR2_X1 XNOR_1_5_N24_PULSESHAPING (.ZN (XNOR_1_5_N24_PULSESHAPING_OUT), .A1 (XNOR_1_4_N24_PULSESHAPING_OUT), .A2 (GND));
       NOR2_X1 XNOR_1_6_N24_PULSESHAPING (.ZN (XNOR_1_6_N24_PULSESHAPING_OUT), .A1 (XNOR_1_5_N24_PULSESHAPING_OUT), .A2 (GND));
       NOR2_X1 XNOR_1_7_N24_PULSESHAPING (.ZN (N24), .A1 (XNOR_1_6_N24_PULSESHAPING_OUT), .A2 (GND));

       wire XNOR_1_1_N27_PULSESHAPING_OUT, XNOR_1_2_N27_PULSESHAPING_OUT, XNOR_1_3_N27_PULSESHAPING_OUT, XNOR_1_4_N27_PULSESHAPING_OUT, XNOR_1_5_N27_PULSESHAPING_OUT, XNOR_1_6_N27_PULSESHAPING_OUT;
       NOR2_X1 XNOR_1_1_N27_PULSESHAPING (.ZN (XNOR_1_1_N27_PULSESHAPING_OUT), .A1 (N27_PWL), .A2 (GND));
       NOR2_X1 XNOR_1_2_N27_PULSESHAPING (.ZN (XNOR_1_2_N27_PULSESHAPING_OUT), .A1 (XNOR_1_1_N27_PULSESHAPING_OUT), .A2 (GND));
       NOR2_X1 XNOR_1_3_N27_PULSESHAPING (.ZN (XNOR_1_3_N27_PULSESHAPING_OUT), .A1 (XNOR_1_2_N27_PULSESHAPING_OUT), .A2 (GND));
       NOR2_X1 XNOR_1_4_N27_PULSESHAPING (.ZN (XNOR_1_4_N27_PULSESHAPING_OUT), .A1 (XNOR_1_3_N27_PULSESHAPING_OUT), .A2 (GND));
       NOR2_X1 XNOR_1_5_N27_PULSESHAPING (.ZN (XNOR_1_5_N27_PULSESHAPING_OUT), .A1 (XNOR_1_4_N27_PULSESHAPING_OUT), .A2 (GND));
       NOR2_X1 XNOR_1_6_N27_PULSESHAPING (.ZN (XNOR_1_6_N27_PULSESHAPING_OUT), .A1 (XNOR_1_5_N27_PULSESHAPING_OUT), .A2 (GND));
       NOR2_X1 XNOR_1_7_N27_PULSESHAPING (.ZN (N27), .A1 (XNOR_1_6_N27_PULSESHAPING_OUT), .A2 (GND));

       wire XNOR_1_1_N30_PULSESHAPING_OUT, XNOR_1_2_N30_PULSESHAPING_OUT, XNOR_1_3_N30_PULSESHAPING_OUT, XNOR_1_4_N30_PULSESHAPING_OUT, XNOR_1_5_N30_PULSESHAPING_OUT, XNOR_1_6_N30_PULSESHAPING_OUT;
       NOR2_X1 XNOR_1_1_N30_PULSESHAPING (.ZN (XNOR_1_1_N30_PULSESHAPING_OUT), .A1 (N30_PWL), .A2 (GND));
       NOR2_X1 XNOR_1_2_N30_PULSESHAPING (.ZN (XNOR_1_2_N30_PULSESHAPING_OUT), .A1 (XNOR_1_1_N30_PULSESHAPING_OUT), .A2 (GND));
       NOR2_X1 XNOR_1_3_N30_PULSESHAPING (.ZN (XNOR_1_3_N30_PULSESHAPING_OUT), .A1 (XNOR_1_2_N30_PULSESHAPING_OUT), .A2 (GND));
       NOR2_X1 XNOR_1_4_N30_PULSESHAPING (.ZN (XNOR_1_4_N30_PULSESHAPING_OUT), .A1 (XNOR_1_3_N30_PULSESHAPING_OUT), .A2 (GND));
       NOR2_X1 XNOR_1_5_N30_PULSESHAPING (.ZN (XNOR_1_5_N30_PULSESHAPING_OUT), .A1 (XNOR_1_4_N30_PULSESHAPING_OUT), .A2 (GND));
       NOR2_X1 XNOR_1_6_N30_PULSESHAPING (.ZN (XNOR_1_6_N30_PULSESHAPING_OUT), .A1 (XNOR_1_5_N30_PULSESHAPING_OUT), .A2 (GND));
       NOR2_X1 XNOR_1_7_N30_PULSESHAPING (.ZN (N30), .A1 (XNOR_1_6_N30_PULSESHAPING_OUT), .A2 (GND));

       wire XNOR_1_1_N34_PULSESHAPING_OUT, XNOR_1_2_N34_PULSESHAPING_OUT, XNOR_1_3_N34_PULSESHAPING_OUT, XNOR_1_4_N34_PULSESHAPING_OUT, XNOR_1_5_N34_PULSESHAPING_OUT, XNOR_1_6_N34_PULSESHAPING_OUT;
       NOR2_X1 XNOR_1_1_N34_PULSESHAPING (.ZN (XNOR_1_1_N34_PULSESHAPING_OUT), .A1 (N34_PWL), .A2 (GND));
       NOR2_X1 XNOR_1_2_N34_PULSESHAPING (.ZN (XNOR_1_2_N34_PULSESHAPING_OUT), .A1 (XNOR_1_1_N34_PULSESHAPING_OUT), .A2 (GND));
       NOR2_X1 XNOR_1_3_N34_PULSESHAPING (.ZN (XNOR_1_3_N34_PULSESHAPING_OUT), .A1 (XNOR_1_2_N34_PULSESHAPING_OUT), .A2 (GND));
       NOR2_X1 XNOR_1_4_N34_PULSESHAPING (.ZN (XNOR_1_4_N34_PULSESHAPING_OUT), .A1 (XNOR_1_3_N34_PULSESHAPING_OUT), .A2 (GND));
       NOR2_X1 XNOR_1_5_N34_PULSESHAPING (.ZN (XNOR_1_5_N34_PULSESHAPING_OUT), .A1 (XNOR_1_4_N34_PULSESHAPING_OUT), .A2 (GND));
       NOR2_X1 XNOR_1_6_N34_PULSESHAPING (.ZN (XNOR_1_6_N34_PULSESHAPING_OUT), .A1 (XNOR_1_5_N34_PULSESHAPING_OUT), .A2 (GND));
       NOR2_X1 XNOR_1_7_N34_PULSESHAPING (.ZN (N34), .A1 (XNOR_1_6_N34_PULSESHAPING_OUT), .A2 (GND));

       wire XNOR_1_1_N37_PULSESHAPING_OUT, XNOR_1_2_N37_PULSESHAPING_OUT, XNOR_1_3_N37_PULSESHAPING_OUT, XNOR_1_4_N37_PULSESHAPING_OUT, XNOR_1_5_N37_PULSESHAPING_OUT, XNOR_1_6_N37_PULSESHAPING_OUT;
       NOR2_X1 XNOR_1_1_N37_PULSESHAPING (.ZN (XNOR_1_1_N37_PULSESHAPING_OUT), .A1 (N37_PWL), .A2 (GND));
       NOR2_X1 XNOR_1_2_N37_PULSESHAPING (.ZN (XNOR_1_2_N37_PULSESHAPING_OUT), .A1 (XNOR_1_1_N37_PULSESHAPING_OUT), .A2 (GND));
       NOR2_X1 XNOR_1_3_N37_PULSESHAPING (.ZN (XNOR_1_3_N37_PULSESHAPING_OUT), .A1 (XNOR_1_2_N37_PULSESHAPING_OUT), .A2 (GND));
       NOR2_X1 XNOR_1_4_N37_PULSESHAPING (.ZN (XNOR_1_4_N37_PULSESHAPING_OUT), .A1 (XNOR_1_3_N37_PULSESHAPING_OUT), .A2 (GND));
       NOR2_X1 XNOR_1_5_N37_PULSESHAPING (.ZN (XNOR_1_5_N37_PULSESHAPING_OUT), .A1 (XNOR_1_4_N37_PULSESHAPING_OUT), .A2 (GND));
       NOR2_X1 XNOR_1_6_N37_PULSESHAPING (.ZN (XNOR_1_6_N37_PULSESHAPING_OUT), .A1 (XNOR_1_5_N37_PULSESHAPING_OUT), .A2 (GND));
       NOR2_X1 XNOR_1_7_N37_PULSESHAPING (.ZN (N37), .A1 (XNOR_1_6_N37_PULSESHAPING_OUT), .A2 (GND));

       wire XNOR_1_1_N40_PULSESHAPING_OUT, XNOR_1_2_N40_PULSESHAPING_OUT, XNOR_1_3_N40_PULSESHAPING_OUT, XNOR_1_4_N40_PULSESHAPING_OUT, XNOR_1_5_N40_PULSESHAPING_OUT, XNOR_1_6_N40_PULSESHAPING_OUT;
       NOR2_X1 XNOR_1_1_N40_PULSESHAPING (.ZN (XNOR_1_1_N40_PULSESHAPING_OUT), .A1 (N40_PWL), .A2 (GND));
       NOR2_X1 XNOR_1_2_N40_PULSESHAPING (.ZN (XNOR_1_2_N40_PULSESHAPING_OUT), .A1 (XNOR_1_1_N40_PULSESHAPING_OUT), .A2 (GND));
       NOR2_X1 XNOR_1_3_N40_PULSESHAPING (.ZN (XNOR_1_3_N40_PULSESHAPING_OUT), .A1 (XNOR_1_2_N40_PULSESHAPING_OUT), .A2 (GND));
       NOR2_X1 XNOR_1_4_N40_PULSESHAPING (.ZN (XNOR_1_4_N40_PULSESHAPING_OUT), .A1 (XNOR_1_3_N40_PULSESHAPING_OUT), .A2 (GND));
       NOR2_X1 XNOR_1_5_N40_PULSESHAPING (.ZN (XNOR_1_5_N40_PULSESHAPING_OUT), .A1 (XNOR_1_4_N40_PULSESHAPING_OUT), .A2 (GND));
       NOR2_X1 XNOR_1_6_N40_PULSESHAPING (.ZN (XNOR_1_6_N40_PULSESHAPING_OUT), .A1 (XNOR_1_5_N40_PULSESHAPING_OUT), .A2 (GND));
       NOR2_X1 XNOR_1_7_N40_PULSESHAPING (.ZN (N40), .A1 (XNOR_1_6_N40_PULSESHAPING_OUT), .A2 (GND));

       wire XNOR_1_1_N43_PULSESHAPING_OUT, XNOR_1_2_N43_PULSESHAPING_OUT, XNOR_1_3_N43_PULSESHAPING_OUT, XNOR_1_4_N43_PULSESHAPING_OUT, XNOR_1_5_N43_PULSESHAPING_OUT, XNOR_1_6_N43_PULSESHAPING_OUT;
       NOR2_X1 XNOR_1_1_N43_PULSESHAPING (.ZN (XNOR_1_1_N43_PULSESHAPING_OUT), .A1 (N43_PWL), .A2 (GND));
       NOR2_X1 XNOR_1_2_N43_PULSESHAPING (.ZN (XNOR_1_2_N43_PULSESHAPING_OUT), .A1 (XNOR_1_1_N43_PULSESHAPING_OUT), .A2 (GND));
       NOR2_X1 XNOR_1_3_N43_PULSESHAPING (.ZN (XNOR_1_3_N43_PULSESHAPING_OUT), .A1 (XNOR_1_2_N43_PULSESHAPING_OUT), .A2 (GND));
       NOR2_X1 XNOR_1_4_N43_PULSESHAPING (.ZN (XNOR_1_4_N43_PULSESHAPING_OUT), .A1 (XNOR_1_3_N43_PULSESHAPING_OUT), .A2 (GND));
       NOR2_X1 XNOR_1_5_N43_PULSESHAPING (.ZN (XNOR_1_5_N43_PULSESHAPING_OUT), .A1 (XNOR_1_4_N43_PULSESHAPING_OUT), .A2 (GND));
       NOR2_X1 XNOR_1_6_N43_PULSESHAPING (.ZN (XNOR_1_6_N43_PULSESHAPING_OUT), .A1 (XNOR_1_5_N43_PULSESHAPING_OUT), .A2 (GND));
       NOR2_X1 XNOR_1_7_N43_PULSESHAPING (.ZN (N43), .A1 (XNOR_1_6_N43_PULSESHAPING_OUT), .A2 (GND));

       wire XNOR_1_1_N47_PULSESHAPING_OUT, XNOR_1_2_N47_PULSESHAPING_OUT, XNOR_1_3_N47_PULSESHAPING_OUT, XNOR_1_4_N47_PULSESHAPING_OUT, XNOR_1_5_N47_PULSESHAPING_OUT, XNOR_1_6_N47_PULSESHAPING_OUT;
       NOR2_X1 XNOR_1_1_N47_PULSESHAPING (.ZN (XNOR_1_1_N47_PULSESHAPING_OUT), .A1 (N47_PWL), .A2 (GND));
       NOR2_X1 XNOR_1_2_N47_PULSESHAPING (.ZN (XNOR_1_2_N47_PULSESHAPING_OUT), .A1 (XNOR_1_1_N47_PULSESHAPING_OUT), .A2 (GND));
       NOR2_X1 XNOR_1_3_N47_PULSESHAPING (.ZN (XNOR_1_3_N47_PULSESHAPING_OUT), .A1 (XNOR_1_2_N47_PULSESHAPING_OUT), .A2 (GND));
       NOR2_X1 XNOR_1_4_N47_PULSESHAPING (.ZN (XNOR_1_4_N47_PULSESHAPING_OUT), .A1 (XNOR_1_3_N47_PULSESHAPING_OUT), .A2 (GND));
       NOR2_X1 XNOR_1_5_N47_PULSESHAPING (.ZN (XNOR_1_5_N47_PULSESHAPING_OUT), .A1 (XNOR_1_4_N47_PULSESHAPING_OUT), .A2 (GND));
       NOR2_X1 XNOR_1_6_N47_PULSESHAPING (.ZN (XNOR_1_6_N47_PULSESHAPING_OUT), .A1 (XNOR_1_5_N47_PULSESHAPING_OUT), .A2 (GND));
       NOR2_X1 XNOR_1_7_N47_PULSESHAPING (.ZN (N47), .A1 (XNOR_1_6_N47_PULSESHAPING_OUT), .A2 (GND));

       wire XNOR_1_1_N50_PULSESHAPING_OUT, XNOR_1_2_N50_PULSESHAPING_OUT, XNOR_1_3_N50_PULSESHAPING_OUT, XNOR_1_4_N50_PULSESHAPING_OUT, XNOR_1_5_N50_PULSESHAPING_OUT, XNOR_1_6_N50_PULSESHAPING_OUT;
       NOR2_X1 XNOR_1_1_N50_PULSESHAPING (.ZN (XNOR_1_1_N50_PULSESHAPING_OUT), .A1 (N50_PWL), .A2 (GND));
       NOR2_X1 XNOR_1_2_N50_PULSESHAPING (.ZN (XNOR_1_2_N50_PULSESHAPING_OUT), .A1 (XNOR_1_1_N50_PULSESHAPING_OUT), .A2 (GND));
       NOR2_X1 XNOR_1_3_N50_PULSESHAPING (.ZN (XNOR_1_3_N50_PULSESHAPING_OUT), .A1 (XNOR_1_2_N50_PULSESHAPING_OUT), .A2 (GND));
       NOR2_X1 XNOR_1_4_N50_PULSESHAPING (.ZN (XNOR_1_4_N50_PULSESHAPING_OUT), .A1 (XNOR_1_3_N50_PULSESHAPING_OUT), .A2 (GND));
       NOR2_X1 XNOR_1_5_N50_PULSESHAPING (.ZN (XNOR_1_5_N50_PULSESHAPING_OUT), .A1 (XNOR_1_4_N50_PULSESHAPING_OUT), .A2 (GND));
       NOR2_X1 XNOR_1_6_N50_PULSESHAPING (.ZN (XNOR_1_6_N50_PULSESHAPING_OUT), .A1 (XNOR_1_5_N50_PULSESHAPING_OUT), .A2 (GND));
       NOR2_X1 XNOR_1_7_N50_PULSESHAPING (.ZN (N50), .A1 (XNOR_1_6_N50_PULSESHAPING_OUT), .A2 (GND));

       wire XNOR_1_1_N53_PULSESHAPING_OUT, XNOR_1_2_N53_PULSESHAPING_OUT, XNOR_1_3_N53_PULSESHAPING_OUT, XNOR_1_4_N53_PULSESHAPING_OUT, XNOR_1_5_N53_PULSESHAPING_OUT, XNOR_1_6_N53_PULSESHAPING_OUT;
       NOR2_X1 XNOR_1_1_N53_PULSESHAPING (.ZN (XNOR_1_1_N53_PULSESHAPING_OUT), .A1 (N53_PWL), .A2 (GND));
       NOR2_X1 XNOR_1_2_N53_PULSESHAPING (.ZN (XNOR_1_2_N53_PULSESHAPING_OUT), .A1 (XNOR_1_1_N53_PULSESHAPING_OUT), .A2 (GND));
       NOR2_X1 XNOR_1_3_N53_PULSESHAPING (.ZN (XNOR_1_3_N53_PULSESHAPING_OUT), .A1 (XNOR_1_2_N53_PULSESHAPING_OUT), .A2 (GND));
       NOR2_X1 XNOR_1_4_N53_PULSESHAPING (.ZN (XNOR_1_4_N53_PULSESHAPING_OUT), .A1 (XNOR_1_3_N53_PULSESHAPING_OUT), .A2 (GND));
       NOR2_X1 XNOR_1_5_N53_PULSESHAPING (.ZN (XNOR_1_5_N53_PULSESHAPING_OUT), .A1 (XNOR_1_4_N53_PULSESHAPING_OUT), .A2 (GND));
       NOR2_X1 XNOR_1_6_N53_PULSESHAPING (.ZN (XNOR_1_6_N53_PULSESHAPING_OUT), .A1 (XNOR_1_5_N53_PULSESHAPING_OUT), .A2 (GND));
       NOR2_X1 XNOR_1_7_N53_PULSESHAPING (.ZN (N53), .A1 (XNOR_1_6_N53_PULSESHAPING_OUT), .A2 (GND));

       wire XNOR_1_1_N56_PULSESHAPING_OUT, XNOR_1_2_N56_PULSESHAPING_OUT, XNOR_1_3_N56_PULSESHAPING_OUT, XNOR_1_4_N56_PULSESHAPING_OUT, XNOR_1_5_N56_PULSESHAPING_OUT, XNOR_1_6_N56_PULSESHAPING_OUT;
       NOR2_X1 XNOR_1_1_N56_PULSESHAPING (.ZN (XNOR_1_1_N56_PULSESHAPING_OUT), .A1 (N56_PWL), .A2 (GND));
       NOR2_X1 XNOR_1_2_N56_PULSESHAPING (.ZN (XNOR_1_2_N56_PULSESHAPING_OUT), .A1 (XNOR_1_1_N56_PULSESHAPING_OUT), .A2 (GND));
       NOR2_X1 XNOR_1_3_N56_PULSESHAPING (.ZN (XNOR_1_3_N56_PULSESHAPING_OUT), .A1 (XNOR_1_2_N56_PULSESHAPING_OUT), .A2 (GND));
       NOR2_X1 XNOR_1_4_N56_PULSESHAPING (.ZN (XNOR_1_4_N56_PULSESHAPING_OUT), .A1 (XNOR_1_3_N56_PULSESHAPING_OUT), .A2 (GND));
       NOR2_X1 XNOR_1_5_N56_PULSESHAPING (.ZN (XNOR_1_5_N56_PULSESHAPING_OUT), .A1 (XNOR_1_4_N56_PULSESHAPING_OUT), .A2 (GND));
       NOR2_X1 XNOR_1_6_N56_PULSESHAPING (.ZN (XNOR_1_6_N56_PULSESHAPING_OUT), .A1 (XNOR_1_5_N56_PULSESHAPING_OUT), .A2 (GND));
       NOR2_X1 XNOR_1_7_N56_PULSESHAPING (.ZN (N56), .A1 (XNOR_1_6_N56_PULSESHAPING_OUT), .A2 (GND));

       wire XNOR_1_1_N60_PULSESHAPING_OUT, XNOR_1_2_N60_PULSESHAPING_OUT, XNOR_1_3_N60_PULSESHAPING_OUT, XNOR_1_4_N60_PULSESHAPING_OUT, XNOR_1_5_N60_PULSESHAPING_OUT, XNOR_1_6_N60_PULSESHAPING_OUT;
       NOR2_X1 XNOR_1_1_N60_PULSESHAPING (.ZN (XNOR_1_1_N60_PULSESHAPING_OUT), .A1 (N60_PWL), .A2 (GND));
       NOR2_X1 XNOR_1_2_N60_PULSESHAPING (.ZN (XNOR_1_2_N60_PULSESHAPING_OUT), .A1 (XNOR_1_1_N60_PULSESHAPING_OUT), .A2 (GND));
       NOR2_X1 XNOR_1_3_N60_PULSESHAPING (.ZN (XNOR_1_3_N60_PULSESHAPING_OUT), .A1 (XNOR_1_2_N60_PULSESHAPING_OUT), .A2 (GND));
       NOR2_X1 XNOR_1_4_N60_PULSESHAPING (.ZN (XNOR_1_4_N60_PULSESHAPING_OUT), .A1 (XNOR_1_3_N60_PULSESHAPING_OUT), .A2 (GND));
       NOR2_X1 XNOR_1_5_N60_PULSESHAPING (.ZN (XNOR_1_5_N60_PULSESHAPING_OUT), .A1 (XNOR_1_4_N60_PULSESHAPING_OUT), .A2 (GND));
       NOR2_X1 XNOR_1_6_N60_PULSESHAPING (.ZN (XNOR_1_6_N60_PULSESHAPING_OUT), .A1 (XNOR_1_5_N60_PULSESHAPING_OUT), .A2 (GND));
       NOR2_X1 XNOR_1_7_N60_PULSESHAPING (.ZN (N60), .A1 (XNOR_1_6_N60_PULSESHAPING_OUT), .A2 (GND));

       wire XNOR_1_1_N63_PULSESHAPING_OUT, XNOR_1_2_N63_PULSESHAPING_OUT, XNOR_1_3_N63_PULSESHAPING_OUT, XNOR_1_4_N63_PULSESHAPING_OUT, XNOR_1_5_N63_PULSESHAPING_OUT, XNOR_1_6_N63_PULSESHAPING_OUT;
       NOR2_X1 XNOR_1_1_N63_PULSESHAPING (.ZN (XNOR_1_1_N63_PULSESHAPING_OUT), .A1 (N63_PWL), .A2 (GND));
       NOR2_X1 XNOR_1_2_N63_PULSESHAPING (.ZN (XNOR_1_2_N63_PULSESHAPING_OUT), .A1 (XNOR_1_1_N63_PULSESHAPING_OUT), .A2 (GND));
       NOR2_X1 XNOR_1_3_N63_PULSESHAPING (.ZN (XNOR_1_3_N63_PULSESHAPING_OUT), .A1 (XNOR_1_2_N63_PULSESHAPING_OUT), .A2 (GND));
       NOR2_X1 XNOR_1_4_N63_PULSESHAPING (.ZN (XNOR_1_4_N63_PULSESHAPING_OUT), .A1 (XNOR_1_3_N63_PULSESHAPING_OUT), .A2 (GND));
       NOR2_X1 XNOR_1_5_N63_PULSESHAPING (.ZN (XNOR_1_5_N63_PULSESHAPING_OUT), .A1 (XNOR_1_4_N63_PULSESHAPING_OUT), .A2 (GND));
       NOR2_X1 XNOR_1_6_N63_PULSESHAPING (.ZN (XNOR_1_6_N63_PULSESHAPING_OUT), .A1 (XNOR_1_5_N63_PULSESHAPING_OUT), .A2 (GND));
       NOR2_X1 XNOR_1_7_N63_PULSESHAPING (.ZN (N63), .A1 (XNOR_1_6_N63_PULSESHAPING_OUT), .A2 (GND));

       wire XNOR_1_1_N66_PULSESHAPING_OUT, XNOR_1_2_N66_PULSESHAPING_OUT, XNOR_1_3_N66_PULSESHAPING_OUT, XNOR_1_4_N66_PULSESHAPING_OUT, XNOR_1_5_N66_PULSESHAPING_OUT, XNOR_1_6_N66_PULSESHAPING_OUT;
       NOR2_X1 XNOR_1_1_N66_PULSESHAPING (.ZN (XNOR_1_1_N66_PULSESHAPING_OUT), .A1 (N66_PWL), .A2 (GND));
       NOR2_X1 XNOR_1_2_N66_PULSESHAPING (.ZN (XNOR_1_2_N66_PULSESHAPING_OUT), .A1 (XNOR_1_1_N66_PULSESHAPING_OUT), .A2 (GND));
       NOR2_X1 XNOR_1_3_N66_PULSESHAPING (.ZN (XNOR_1_3_N66_PULSESHAPING_OUT), .A1 (XNOR_1_2_N66_PULSESHAPING_OUT), .A2 (GND));
       NOR2_X1 XNOR_1_4_N66_PULSESHAPING (.ZN (XNOR_1_4_N66_PULSESHAPING_OUT), .A1 (XNOR_1_3_N66_PULSESHAPING_OUT), .A2 (GND));
       NOR2_X1 XNOR_1_5_N66_PULSESHAPING (.ZN (XNOR_1_5_N66_PULSESHAPING_OUT), .A1 (XNOR_1_4_N66_PULSESHAPING_OUT), .A2 (GND));
       NOR2_X1 XNOR_1_6_N66_PULSESHAPING (.ZN (XNOR_1_6_N66_PULSESHAPING_OUT), .A1 (XNOR_1_5_N66_PULSESHAPING_OUT), .A2 (GND));
       NOR2_X1 XNOR_1_7_N66_PULSESHAPING (.ZN (N66), .A1 (XNOR_1_6_N66_PULSESHAPING_OUT), .A2 (GND));

       wire XNOR_1_1_N69_PULSESHAPING_OUT, XNOR_1_2_N69_PULSESHAPING_OUT, XNOR_1_3_N69_PULSESHAPING_OUT, XNOR_1_4_N69_PULSESHAPING_OUT, XNOR_1_5_N69_PULSESHAPING_OUT, XNOR_1_6_N69_PULSESHAPING_OUT;
       NOR2_X1 XNOR_1_1_N69_PULSESHAPING (.ZN (XNOR_1_1_N69_PULSESHAPING_OUT), .A1 (N69_PWL), .A2 (GND));
       NOR2_X1 XNOR_1_2_N69_PULSESHAPING (.ZN (XNOR_1_2_N69_PULSESHAPING_OUT), .A1 (XNOR_1_1_N69_PULSESHAPING_OUT), .A2 (GND));
       NOR2_X1 XNOR_1_3_N69_PULSESHAPING (.ZN (XNOR_1_3_N69_PULSESHAPING_OUT), .A1 (XNOR_1_2_N69_PULSESHAPING_OUT), .A2 (GND));
       NOR2_X1 XNOR_1_4_N69_PULSESHAPING (.ZN (XNOR_1_4_N69_PULSESHAPING_OUT), .A1 (XNOR_1_3_N69_PULSESHAPING_OUT), .A2 (GND));
       NOR2_X1 XNOR_1_5_N69_PULSESHAPING (.ZN (XNOR_1_5_N69_PULSESHAPING_OUT), .A1 (XNOR_1_4_N69_PULSESHAPING_OUT), .A2 (GND));
       NOR2_X1 XNOR_1_6_N69_PULSESHAPING (.ZN (XNOR_1_6_N69_PULSESHAPING_OUT), .A1 (XNOR_1_5_N69_PULSESHAPING_OUT), .A2 (GND));
       NOR2_X1 XNOR_1_7_N69_PULSESHAPING (.ZN (N69), .A1 (XNOR_1_6_N69_PULSESHAPING_OUT), .A2 (GND));

       wire XNOR_1_1_N73_PULSESHAPING_OUT, XNOR_1_2_N73_PULSESHAPING_OUT, XNOR_1_3_N73_PULSESHAPING_OUT, XNOR_1_4_N73_PULSESHAPING_OUT, XNOR_1_5_N73_PULSESHAPING_OUT, XNOR_1_6_N73_PULSESHAPING_OUT;
       NOR2_X1 XNOR_1_1_N73_PULSESHAPING (.ZN (XNOR_1_1_N73_PULSESHAPING_OUT), .A1 (N73_PWL), .A2 (GND));
       NOR2_X1 XNOR_1_2_N73_PULSESHAPING (.ZN (XNOR_1_2_N73_PULSESHAPING_OUT), .A1 (XNOR_1_1_N73_PULSESHAPING_OUT), .A2 (GND));
       NOR2_X1 XNOR_1_3_N73_PULSESHAPING (.ZN (XNOR_1_3_N73_PULSESHAPING_OUT), .A1 (XNOR_1_2_N73_PULSESHAPING_OUT), .A2 (GND));
       NOR2_X1 XNOR_1_4_N73_PULSESHAPING (.ZN (XNOR_1_4_N73_PULSESHAPING_OUT), .A1 (XNOR_1_3_N73_PULSESHAPING_OUT), .A2 (GND));
       NOR2_X1 XNOR_1_5_N73_PULSESHAPING (.ZN (XNOR_1_5_N73_PULSESHAPING_OUT), .A1 (XNOR_1_4_N73_PULSESHAPING_OUT), .A2 (GND));
       NOR2_X1 XNOR_1_6_N73_PULSESHAPING (.ZN (XNOR_1_6_N73_PULSESHAPING_OUT), .A1 (XNOR_1_5_N73_PULSESHAPING_OUT), .A2 (GND));
       NOR2_X1 XNOR_1_7_N73_PULSESHAPING (.ZN (N73), .A1 (XNOR_1_6_N73_PULSESHAPING_OUT), .A2 (GND));

       wire XNOR_1_1_N76_PULSESHAPING_OUT, XNOR_1_2_N76_PULSESHAPING_OUT, XNOR_1_3_N76_PULSESHAPING_OUT, XNOR_1_4_N76_PULSESHAPING_OUT, XNOR_1_5_N76_PULSESHAPING_OUT, XNOR_1_6_N76_PULSESHAPING_OUT;
       NOR2_X1 XNOR_1_1_N76_PULSESHAPING (.ZN (XNOR_1_1_N76_PULSESHAPING_OUT), .A1 (N76_PWL), .A2 (GND));
       NOR2_X1 XNOR_1_2_N76_PULSESHAPING (.ZN (XNOR_1_2_N76_PULSESHAPING_OUT), .A1 (XNOR_1_1_N76_PULSESHAPING_OUT), .A2 (GND));
       NOR2_X1 XNOR_1_3_N76_PULSESHAPING (.ZN (XNOR_1_3_N76_PULSESHAPING_OUT), .A1 (XNOR_1_2_N76_PULSESHAPING_OUT), .A2 (GND));
       NOR2_X1 XNOR_1_4_N76_PULSESHAPING (.ZN (XNOR_1_4_N76_PULSESHAPING_OUT), .A1 (XNOR_1_3_N76_PULSESHAPING_OUT), .A2 (GND));
       NOR2_X1 XNOR_1_5_N76_PULSESHAPING (.ZN (XNOR_1_5_N76_PULSESHAPING_OUT), .A1 (XNOR_1_4_N76_PULSESHAPING_OUT), .A2 (GND));
       NOR2_X1 XNOR_1_6_N76_PULSESHAPING (.ZN (XNOR_1_6_N76_PULSESHAPING_OUT), .A1 (XNOR_1_5_N76_PULSESHAPING_OUT), .A2 (GND));
       NOR2_X1 XNOR_1_7_N76_PULSESHAPING (.ZN (N76), .A1 (XNOR_1_6_N76_PULSESHAPING_OUT), .A2 (GND));

       wire XNOR_1_1_N79_PULSESHAPING_OUT, XNOR_1_2_N79_PULSESHAPING_OUT, XNOR_1_3_N79_PULSESHAPING_OUT, XNOR_1_4_N79_PULSESHAPING_OUT, XNOR_1_5_N79_PULSESHAPING_OUT, XNOR_1_6_N79_PULSESHAPING_OUT;
       NOR2_X1 XNOR_1_1_N79_PULSESHAPING (.ZN (XNOR_1_1_N79_PULSESHAPING_OUT), .A1 (N79_PWL), .A2 (GND));
       NOR2_X1 XNOR_1_2_N79_PULSESHAPING (.ZN (XNOR_1_2_N79_PULSESHAPING_OUT), .A1 (XNOR_1_1_N79_PULSESHAPING_OUT), .A2 (GND));
       NOR2_X1 XNOR_1_3_N79_PULSESHAPING (.ZN (XNOR_1_3_N79_PULSESHAPING_OUT), .A1 (XNOR_1_2_N79_PULSESHAPING_OUT), .A2 (GND));
       NOR2_X1 XNOR_1_4_N79_PULSESHAPING (.ZN (XNOR_1_4_N79_PULSESHAPING_OUT), .A1 (XNOR_1_3_N79_PULSESHAPING_OUT), .A2 (GND));
       NOR2_X1 XNOR_1_5_N79_PULSESHAPING (.ZN (XNOR_1_5_N79_PULSESHAPING_OUT), .A1 (XNOR_1_4_N79_PULSESHAPING_OUT), .A2 (GND));
       NOR2_X1 XNOR_1_6_N79_PULSESHAPING (.ZN (XNOR_1_6_N79_PULSESHAPING_OUT), .A1 (XNOR_1_5_N79_PULSESHAPING_OUT), .A2 (GND));
       NOR2_X1 XNOR_1_7_N79_PULSESHAPING (.ZN (N79), .A1 (XNOR_1_6_N79_PULSESHAPING_OUT), .A2 (GND));

       wire XNOR_1_1_N82_PULSESHAPING_OUT, XNOR_1_2_N82_PULSESHAPING_OUT, XNOR_1_3_N82_PULSESHAPING_OUT, XNOR_1_4_N82_PULSESHAPING_OUT, XNOR_1_5_N82_PULSESHAPING_OUT, XNOR_1_6_N82_PULSESHAPING_OUT;
       NOR2_X1 XNOR_1_1_N82_PULSESHAPING (.ZN (XNOR_1_1_N82_PULSESHAPING_OUT), .A1 (N82_PWL), .A2 (GND));
       NOR2_X1 XNOR_1_2_N82_PULSESHAPING (.ZN (XNOR_1_2_N82_PULSESHAPING_OUT), .A1 (XNOR_1_1_N82_PULSESHAPING_OUT), .A2 (GND));
       NOR2_X1 XNOR_1_3_N82_PULSESHAPING (.ZN (XNOR_1_3_N82_PULSESHAPING_OUT), .A1 (XNOR_1_2_N82_PULSESHAPING_OUT), .A2 (GND));
       NOR2_X1 XNOR_1_4_N82_PULSESHAPING (.ZN (XNOR_1_4_N82_PULSESHAPING_OUT), .A1 (XNOR_1_3_N82_PULSESHAPING_OUT), .A2 (GND));
       NOR2_X1 XNOR_1_5_N82_PULSESHAPING (.ZN (XNOR_1_5_N82_PULSESHAPING_OUT), .A1 (XNOR_1_4_N82_PULSESHAPING_OUT), .A2 (GND));
       NOR2_X1 XNOR_1_6_N82_PULSESHAPING (.ZN (XNOR_1_6_N82_PULSESHAPING_OUT), .A1 (XNOR_1_5_N82_PULSESHAPING_OUT), .A2 (GND));
       NOR2_X1 XNOR_1_7_N82_PULSESHAPING (.ZN (N82), .A1 (XNOR_1_6_N82_PULSESHAPING_OUT), .A2 (GND));

       wire XNOR_1_1_N86_PULSESHAPING_OUT, XNOR_1_2_N86_PULSESHAPING_OUT, XNOR_1_3_N86_PULSESHAPING_OUT, XNOR_1_4_N86_PULSESHAPING_OUT, XNOR_1_5_N86_PULSESHAPING_OUT, XNOR_1_6_N86_PULSESHAPING_OUT;
       NOR2_X1 XNOR_1_1_N86_PULSESHAPING (.ZN (XNOR_1_1_N86_PULSESHAPING_OUT), .A1 (N86_PWL), .A2 (GND));
       NOR2_X1 XNOR_1_2_N86_PULSESHAPING (.ZN (XNOR_1_2_N86_PULSESHAPING_OUT), .A1 (XNOR_1_1_N86_PULSESHAPING_OUT), .A2 (GND));
       NOR2_X1 XNOR_1_3_N86_PULSESHAPING (.ZN (XNOR_1_3_N86_PULSESHAPING_OUT), .A1 (XNOR_1_2_N86_PULSESHAPING_OUT), .A2 (GND));
       NOR2_X1 XNOR_1_4_N86_PULSESHAPING (.ZN (XNOR_1_4_N86_PULSESHAPING_OUT), .A1 (XNOR_1_3_N86_PULSESHAPING_OUT), .A2 (GND));
       NOR2_X1 XNOR_1_5_N86_PULSESHAPING (.ZN (XNOR_1_5_N86_PULSESHAPING_OUT), .A1 (XNOR_1_4_N86_PULSESHAPING_OUT), .A2 (GND));
       NOR2_X1 XNOR_1_6_N86_PULSESHAPING (.ZN (XNOR_1_6_N86_PULSESHAPING_OUT), .A1 (XNOR_1_5_N86_PULSESHAPING_OUT), .A2 (GND));
       NOR2_X1 XNOR_1_7_N86_PULSESHAPING (.ZN (N86), .A1 (XNOR_1_6_N86_PULSESHAPING_OUT), .A2 (GND));

       wire XNOR_1_1_N89_PULSESHAPING_OUT, XNOR_1_2_N89_PULSESHAPING_OUT, XNOR_1_3_N89_PULSESHAPING_OUT, XNOR_1_4_N89_PULSESHAPING_OUT, XNOR_1_5_N89_PULSESHAPING_OUT, XNOR_1_6_N89_PULSESHAPING_OUT;
       NOR2_X1 XNOR_1_1_N89_PULSESHAPING (.ZN (XNOR_1_1_N89_PULSESHAPING_OUT), .A1 (N89_PWL), .A2 (GND));
       NOR2_X1 XNOR_1_2_N89_PULSESHAPING (.ZN (XNOR_1_2_N89_PULSESHAPING_OUT), .A1 (XNOR_1_1_N89_PULSESHAPING_OUT), .A2 (GND));
       NOR2_X1 XNOR_1_3_N89_PULSESHAPING (.ZN (XNOR_1_3_N89_PULSESHAPING_OUT), .A1 (XNOR_1_2_N89_PULSESHAPING_OUT), .A2 (GND));
       NOR2_X1 XNOR_1_4_N89_PULSESHAPING (.ZN (XNOR_1_4_N89_PULSESHAPING_OUT), .A1 (XNOR_1_3_N89_PULSESHAPING_OUT), .A2 (GND));
       NOR2_X1 XNOR_1_5_N89_PULSESHAPING (.ZN (XNOR_1_5_N89_PULSESHAPING_OUT), .A1 (XNOR_1_4_N89_PULSESHAPING_OUT), .A2 (GND));
       NOR2_X1 XNOR_1_6_N89_PULSESHAPING (.ZN (XNOR_1_6_N89_PULSESHAPING_OUT), .A1 (XNOR_1_5_N89_PULSESHAPING_OUT), .A2 (GND));
       NOR2_X1 XNOR_1_7_N89_PULSESHAPING (.ZN (N89), .A1 (XNOR_1_6_N89_PULSESHAPING_OUT), .A2 (GND));

       wire XNOR_1_1_N92_PULSESHAPING_OUT, XNOR_1_2_N92_PULSESHAPING_OUT, XNOR_1_3_N92_PULSESHAPING_OUT, XNOR_1_4_N92_PULSESHAPING_OUT, XNOR_1_5_N92_PULSESHAPING_OUT, XNOR_1_6_N92_PULSESHAPING_OUT;
       NOR2_X1 XNOR_1_1_N92_PULSESHAPING (.ZN (XNOR_1_1_N92_PULSESHAPING_OUT), .A1 (N92_PWL), .A2 (GND));
       NOR2_X1 XNOR_1_2_N92_PULSESHAPING (.ZN (XNOR_1_2_N92_PULSESHAPING_OUT), .A1 (XNOR_1_1_N92_PULSESHAPING_OUT), .A2 (GND));
       NOR2_X1 XNOR_1_3_N92_PULSESHAPING (.ZN (XNOR_1_3_N92_PULSESHAPING_OUT), .A1 (XNOR_1_2_N92_PULSESHAPING_OUT), .A2 (GND));
       NOR2_X1 XNOR_1_4_N92_PULSESHAPING (.ZN (XNOR_1_4_N92_PULSESHAPING_OUT), .A1 (XNOR_1_3_N92_PULSESHAPING_OUT), .A2 (GND));
       NOR2_X1 XNOR_1_5_N92_PULSESHAPING (.ZN (XNOR_1_5_N92_PULSESHAPING_OUT), .A1 (XNOR_1_4_N92_PULSESHAPING_OUT), .A2 (GND));
       NOR2_X1 XNOR_1_6_N92_PULSESHAPING (.ZN (XNOR_1_6_N92_PULSESHAPING_OUT), .A1 (XNOR_1_5_N92_PULSESHAPING_OUT), .A2 (GND));
       NOR2_X1 XNOR_1_7_N92_PULSESHAPING (.ZN (N92), .A1 (XNOR_1_6_N92_PULSESHAPING_OUT), .A2 (GND));

       wire XNOR_1_1_N95_PULSESHAPING_OUT, XNOR_1_2_N95_PULSESHAPING_OUT, XNOR_1_3_N95_PULSESHAPING_OUT, XNOR_1_4_N95_PULSESHAPING_OUT, XNOR_1_5_N95_PULSESHAPING_OUT, XNOR_1_6_N95_PULSESHAPING_OUT;
       NOR2_X1 XNOR_1_1_N95_PULSESHAPING (.ZN (XNOR_1_1_N95_PULSESHAPING_OUT), .A1 (N95_PWL), .A2 (GND));
       NOR2_X1 XNOR_1_2_N95_PULSESHAPING (.ZN (XNOR_1_2_N95_PULSESHAPING_OUT), .A1 (XNOR_1_1_N95_PULSESHAPING_OUT), .A2 (GND));
       NOR2_X1 XNOR_1_3_N95_PULSESHAPING (.ZN (XNOR_1_3_N95_PULSESHAPING_OUT), .A1 (XNOR_1_2_N95_PULSESHAPING_OUT), .A2 (GND));
       NOR2_X1 XNOR_1_4_N95_PULSESHAPING (.ZN (XNOR_1_4_N95_PULSESHAPING_OUT), .A1 (XNOR_1_3_N95_PULSESHAPING_OUT), .A2 (GND));
       NOR2_X1 XNOR_1_5_N95_PULSESHAPING (.ZN (XNOR_1_5_N95_PULSESHAPING_OUT), .A1 (XNOR_1_4_N95_PULSESHAPING_OUT), .A2 (GND));
       NOR2_X1 XNOR_1_6_N95_PULSESHAPING (.ZN (XNOR_1_6_N95_PULSESHAPING_OUT), .A1 (XNOR_1_5_N95_PULSESHAPING_OUT), .A2 (GND));
       NOR2_X1 XNOR_1_7_N95_PULSESHAPING (.ZN (N95), .A1 (XNOR_1_6_N95_PULSESHAPING_OUT), .A2 (GND));

       wire XNOR_1_1_N99_PULSESHAPING_OUT, XNOR_1_2_N99_PULSESHAPING_OUT, XNOR_1_3_N99_PULSESHAPING_OUT, XNOR_1_4_N99_PULSESHAPING_OUT, XNOR_1_5_N99_PULSESHAPING_OUT, XNOR_1_6_N99_PULSESHAPING_OUT;
       NOR2_X1 XNOR_1_1_N99_PULSESHAPING (.ZN (XNOR_1_1_N99_PULSESHAPING_OUT), .A1 (N99_PWL), .A2 (GND));
       NOR2_X1 XNOR_1_2_N99_PULSESHAPING (.ZN (XNOR_1_2_N99_PULSESHAPING_OUT), .A1 (XNOR_1_1_N99_PULSESHAPING_OUT), .A2 (GND));
       NOR2_X1 XNOR_1_3_N99_PULSESHAPING (.ZN (XNOR_1_3_N99_PULSESHAPING_OUT), .A1 (XNOR_1_2_N99_PULSESHAPING_OUT), .A2 (GND));
       NOR2_X1 XNOR_1_4_N99_PULSESHAPING (.ZN (XNOR_1_4_N99_PULSESHAPING_OUT), .A1 (XNOR_1_3_N99_PULSESHAPING_OUT), .A2 (GND));
       NOR2_X1 XNOR_1_5_N99_PULSESHAPING (.ZN (XNOR_1_5_N99_PULSESHAPING_OUT), .A1 (XNOR_1_4_N99_PULSESHAPING_OUT), .A2 (GND));
       NOR2_X1 XNOR_1_6_N99_PULSESHAPING (.ZN (XNOR_1_6_N99_PULSESHAPING_OUT), .A1 (XNOR_1_5_N99_PULSESHAPING_OUT), .A2 (GND));
       NOR2_X1 XNOR_1_7_N99_PULSESHAPING (.ZN (N99), .A1 (XNOR_1_6_N99_PULSESHAPING_OUT), .A2 (GND));

       wire XNOR_1_1_N102_PULSESHAPING_OUT, XNOR_1_2_N102_PULSESHAPING_OUT, XNOR_1_3_N102_PULSESHAPING_OUT, XNOR_1_4_N102_PULSESHAPING_OUT, XNOR_1_5_N102_PULSESHAPING_OUT, XNOR_1_6_N102_PULSESHAPING_OUT;
       NOR2_X1 XNOR_1_1_N102_PULSESHAPING (.ZN (XNOR_1_1_N102_PULSESHAPING_OUT), .A1 (N102_PWL), .A2 (GND));
       NOR2_X1 XNOR_1_2_N102_PULSESHAPING (.ZN (XNOR_1_2_N102_PULSESHAPING_OUT), .A1 (XNOR_1_1_N102_PULSESHAPING_OUT), .A2 (GND));
       NOR2_X1 XNOR_1_3_N102_PULSESHAPING (.ZN (XNOR_1_3_N102_PULSESHAPING_OUT), .A1 (XNOR_1_2_N102_PULSESHAPING_OUT), .A2 (GND));
       NOR2_X1 XNOR_1_4_N102_PULSESHAPING (.ZN (XNOR_1_4_N102_PULSESHAPING_OUT), .A1 (XNOR_1_3_N102_PULSESHAPING_OUT), .A2 (GND));
       NOR2_X1 XNOR_1_5_N102_PULSESHAPING (.ZN (XNOR_1_5_N102_PULSESHAPING_OUT), .A1 (XNOR_1_4_N102_PULSESHAPING_OUT), .A2 (GND));
       NOR2_X1 XNOR_1_6_N102_PULSESHAPING (.ZN (XNOR_1_6_N102_PULSESHAPING_OUT), .A1 (XNOR_1_5_N102_PULSESHAPING_OUT), .A2 (GND));
       NOR2_X1 XNOR_1_7_N102_PULSESHAPING (.ZN (N102), .A1 (XNOR_1_6_N102_PULSESHAPING_OUT), .A2 (GND));

       wire XNOR_1_1_N105_PULSESHAPING_OUT, XNOR_1_2_N105_PULSESHAPING_OUT, XNOR_1_3_N105_PULSESHAPING_OUT, XNOR_1_4_N105_PULSESHAPING_OUT, XNOR_1_5_N105_PULSESHAPING_OUT, XNOR_1_6_N105_PULSESHAPING_OUT;
       NOR2_X1 XNOR_1_1_N105_PULSESHAPING (.ZN (XNOR_1_1_N105_PULSESHAPING_OUT), .A1 (N105_PWL), .A2 (GND));
       NOR2_X1 XNOR_1_2_N105_PULSESHAPING (.ZN (XNOR_1_2_N105_PULSESHAPING_OUT), .A1 (XNOR_1_1_N105_PULSESHAPING_OUT), .A2 (GND));
       NOR2_X1 XNOR_1_3_N105_PULSESHAPING (.ZN (XNOR_1_3_N105_PULSESHAPING_OUT), .A1 (XNOR_1_2_N105_PULSESHAPING_OUT), .A2 (GND));
       NOR2_X1 XNOR_1_4_N105_PULSESHAPING (.ZN (XNOR_1_4_N105_PULSESHAPING_OUT), .A1 (XNOR_1_3_N105_PULSESHAPING_OUT), .A2 (GND));
       NOR2_X1 XNOR_1_5_N105_PULSESHAPING (.ZN (XNOR_1_5_N105_PULSESHAPING_OUT), .A1 (XNOR_1_4_N105_PULSESHAPING_OUT), .A2 (GND));
       NOR2_X1 XNOR_1_6_N105_PULSESHAPING (.ZN (XNOR_1_6_N105_PULSESHAPING_OUT), .A1 (XNOR_1_5_N105_PULSESHAPING_OUT), .A2 (GND));
       NOR2_X1 XNOR_1_7_N105_PULSESHAPING (.ZN (N105), .A1 (XNOR_1_6_N105_PULSESHAPING_OUT), .A2 (GND));

       wire XNOR_1_1_N108_PULSESHAPING_OUT, XNOR_1_2_N108_PULSESHAPING_OUT, XNOR_1_3_N108_PULSESHAPING_OUT, XNOR_1_4_N108_PULSESHAPING_OUT, XNOR_1_5_N108_PULSESHAPING_OUT, XNOR_1_6_N108_PULSESHAPING_OUT;
       NOR2_X1 XNOR_1_1_N108_PULSESHAPING (.ZN (XNOR_1_1_N108_PULSESHAPING_OUT), .A1 (N108_PWL), .A2 (GND));
       NOR2_X1 XNOR_1_2_N108_PULSESHAPING (.ZN (XNOR_1_2_N108_PULSESHAPING_OUT), .A1 (XNOR_1_1_N108_PULSESHAPING_OUT), .A2 (GND));
       NOR2_X1 XNOR_1_3_N108_PULSESHAPING (.ZN (XNOR_1_3_N108_PULSESHAPING_OUT), .A1 (XNOR_1_2_N108_PULSESHAPING_OUT), .A2 (GND));
       NOR2_X1 XNOR_1_4_N108_PULSESHAPING (.ZN (XNOR_1_4_N108_PULSESHAPING_OUT), .A1 (XNOR_1_3_N108_PULSESHAPING_OUT), .A2 (GND));
       NOR2_X1 XNOR_1_5_N108_PULSESHAPING (.ZN (XNOR_1_5_N108_PULSESHAPING_OUT), .A1 (XNOR_1_4_N108_PULSESHAPING_OUT), .A2 (GND));
       NOR2_X1 XNOR_1_6_N108_PULSESHAPING (.ZN (XNOR_1_6_N108_PULSESHAPING_OUT), .A1 (XNOR_1_5_N108_PULSESHAPING_OUT), .A2 (GND));
       NOR2_X1 XNOR_1_7_N108_PULSESHAPING (.ZN (N108), .A1 (XNOR_1_6_N108_PULSESHAPING_OUT), .A2 (GND));

       wire XNOR_1_1_N112_PULSESHAPING_OUT, XNOR_1_2_N112_PULSESHAPING_OUT, XNOR_1_3_N112_PULSESHAPING_OUT, XNOR_1_4_N112_PULSESHAPING_OUT, XNOR_1_5_N112_PULSESHAPING_OUT, XNOR_1_6_N112_PULSESHAPING_OUT;
       NOR2_X1 XNOR_1_1_N112_PULSESHAPING (.ZN (XNOR_1_1_N112_PULSESHAPING_OUT), .A1 (N112_PWL), .A2 (GND));
       NOR2_X1 XNOR_1_2_N112_PULSESHAPING (.ZN (XNOR_1_2_N112_PULSESHAPING_OUT), .A1 (XNOR_1_1_N112_PULSESHAPING_OUT), .A2 (GND));
       NOR2_X1 XNOR_1_3_N112_PULSESHAPING (.ZN (XNOR_1_3_N112_PULSESHAPING_OUT), .A1 (XNOR_1_2_N112_PULSESHAPING_OUT), .A2 (GND));
       NOR2_X1 XNOR_1_4_N112_PULSESHAPING (.ZN (XNOR_1_4_N112_PULSESHAPING_OUT), .A1 (XNOR_1_3_N112_PULSESHAPING_OUT), .A2 (GND));
       NOR2_X1 XNOR_1_5_N112_PULSESHAPING (.ZN (XNOR_1_5_N112_PULSESHAPING_OUT), .A1 (XNOR_1_4_N112_PULSESHAPING_OUT), .A2 (GND));
       NOR2_X1 XNOR_1_6_N112_PULSESHAPING (.ZN (XNOR_1_6_N112_PULSESHAPING_OUT), .A1 (XNOR_1_5_N112_PULSESHAPING_OUT), .A2 (GND));
       NOR2_X1 XNOR_1_7_N112_PULSESHAPING (.ZN (N112), .A1 (XNOR_1_6_N112_PULSESHAPING_OUT), .A2 (GND));

       wire XNOR_1_1_N115_PULSESHAPING_OUT, XNOR_1_2_N115_PULSESHAPING_OUT, XNOR_1_3_N115_PULSESHAPING_OUT, XNOR_1_4_N115_PULSESHAPING_OUT, XNOR_1_5_N115_PULSESHAPING_OUT, XNOR_1_6_N115_PULSESHAPING_OUT;
       NOR2_X1 XNOR_1_1_N115_PULSESHAPING (.ZN (XNOR_1_1_N115_PULSESHAPING_OUT), .A1 (N115_PWL), .A2 (GND));
       NOR2_X1 XNOR_1_2_N115_PULSESHAPING (.ZN (XNOR_1_2_N115_PULSESHAPING_OUT), .A1 (XNOR_1_1_N115_PULSESHAPING_OUT), .A2 (GND));
       NOR2_X1 XNOR_1_3_N115_PULSESHAPING (.ZN (XNOR_1_3_N115_PULSESHAPING_OUT), .A1 (XNOR_1_2_N115_PULSESHAPING_OUT), .A2 (GND));
       NOR2_X1 XNOR_1_4_N115_PULSESHAPING (.ZN (XNOR_1_4_N115_PULSESHAPING_OUT), .A1 (XNOR_1_3_N115_PULSESHAPING_OUT), .A2 (GND));
       NOR2_X1 XNOR_1_5_N115_PULSESHAPING (.ZN (XNOR_1_5_N115_PULSESHAPING_OUT), .A1 (XNOR_1_4_N115_PULSESHAPING_OUT), .A2 (GND));
       NOR2_X1 XNOR_1_6_N115_PULSESHAPING (.ZN (XNOR_1_6_N115_PULSESHAPING_OUT), .A1 (XNOR_1_5_N115_PULSESHAPING_OUT), .A2 (GND));
       NOR2_X1 XNOR_1_7_N115_PULSESHAPING (.ZN (N115), .A1 (XNOR_1_6_N115_PULSESHAPING_OUT), .A2 (GND));



       NOR2_X1 XNOR_NUM1 (.ZN (N118), .A1 (N1), .A2 (GND));
       NOR2_X1 XNOR_NUM2 (.ZN (N119), .A1 (N4), .A2 (GND));
       NOR2_X1 XNOR_NUM3 (.ZN (N122), .A1 (N11), .A2 (GND));
       NOR2_X1 XNOR_NUM4 (.ZN (N123), .A1 (N17), .A2 (GND));
       NOR2_X1 XNOR_NUM5 (.ZN (N126), .A1 (N24), .A2 (GND));
       NOR2_X1 XNOR_NUM6 (.ZN (N127), .A1 (N30), .A2 (GND));
       NOR2_X1 XNOR_NUM7 (.ZN (N130), .A1 (N37), .A2 (GND));
       NOR2_X1 XNOR_NUM8 (.ZN (N131), .A1 (N43), .A2 (GND));
       NOR2_X1 XNOR_NUM9 (.ZN (N134), .A1 (N50), .A2 (GND));
       NOR2_X1 XNOR_NUM10 (.ZN (N135), .A1 (N56), .A2 (GND));
       NOR2_X1 XNOR_NUM11 (.ZN (N138), .A1 (N63), .A2 (GND));
       NOR2_X1 XNOR_NUM12 (.ZN (N139), .A1 (N69), .A2 (GND));
       NOR2_X1 XNOR_NUM13 (.ZN (N142), .A1 (N76), .A2 (GND));
       NOR2_X1 XNOR_NUM14 (.ZN (N143), .A1 (N82), .A2 (GND));
       NOR2_X1 XNOR_NUM15 (.ZN (N146), .A1 (N89), .A2 (GND));
       NOR2_X1 XNOR_NUM16 (.ZN (N147), .A1 (N95), .A2 (GND));
       NOR2_X1 XNOR_NUM17 (.ZN (N150), .A1 (N102), .A2 (GND));
       NOR2_X1 XNOR_NUM18 (.ZN (N151), .A1 (N108), .A2 (GND));
       wire XNOR_1_1_NUM19_OUT, XNOR_1_2_NUM19_OUT, XNOR_1_3_NUM19_OUT;
       NOR2_X1 XNOR_1_1_NUM19 (.ZN (XNOR_1_1_NUM19_OUT), .A1 (N118), .A2 (GND));
       NOR2_X1 XNOR_1_2_NUM19 (.ZN (XNOR_1_2_NUM19_OUT), .A1 (GND), .A2 (N4));
       NOR2_X1 XNOR_1_3_NUM19 (.ZN (XNOR_1_3_NUM19_OUT), .A1 (XNOR_1_1_NUM19_OUT), .A2 (XNOR_1_2_NUM19_OUT));
       NOR2_X1 XNOR_1_4_NUM19 (.ZN (N154), .A1 (XNOR_1_3_NUM19_OUT), .A2 (GND));
       NOR2_X1 XNOR_NUM20 (.ZN (N157), .A1 (N8), .A2 (N119));
       NOR2_X1 XNOR_NUM21 (.ZN (N158), .A1 (N14), .A2 (N119));
       wire XNOR_1_1_NUM22_OUT, XNOR_1_2_NUM22_OUT, XNOR_1_3_NUM22_OUT;
       NOR2_X1 XNOR_1_1_NUM22 (.ZN (XNOR_1_1_NUM22_OUT), .A1 (N122), .A2 (GND));
       NOR2_X1 XNOR_1_2_NUM22 (.ZN (XNOR_1_2_NUM22_OUT), .A1 (GND), .A2 (N17));
       NOR2_X1 XNOR_1_3_NUM22 (.ZN (XNOR_1_3_NUM22_OUT), .A1 (XNOR_1_1_NUM22_OUT), .A2 (XNOR_1_2_NUM22_OUT));
       NOR2_X1 XNOR_1_4_NUM22 (.ZN (N159), .A1 (XNOR_1_3_NUM22_OUT), .A2 (GND));
       wire XNOR_1_1_NUM23_OUT, XNOR_1_2_NUM23_OUT, XNOR_1_3_NUM23_OUT;
       NOR2_X1 XNOR_1_1_NUM23 (.ZN (XNOR_1_1_NUM23_OUT), .A1 (N126), .A2 (GND));
       NOR2_X1 XNOR_1_2_NUM23 (.ZN (XNOR_1_2_NUM23_OUT), .A1 (GND), .A2 (N30));
       NOR2_X1 XNOR_1_3_NUM23 (.ZN (XNOR_1_3_NUM23_OUT), .A1 (XNOR_1_1_NUM23_OUT), .A2 (XNOR_1_2_NUM23_OUT));
       NOR2_X1 XNOR_1_4_NUM23 (.ZN (N162), .A1 (XNOR_1_3_NUM23_OUT), .A2 (GND));
       wire XNOR_1_1_NUM24_OUT, XNOR_1_2_NUM24_OUT, XNOR_1_3_NUM24_OUT;
       NOR2_X1 XNOR_1_1_NUM24 (.ZN (XNOR_1_1_NUM24_OUT), .A1 (N130), .A2 (GND));
       NOR2_X1 XNOR_1_2_NUM24 (.ZN (XNOR_1_2_NUM24_OUT), .A1 (GND), .A2 (N43));
       NOR2_X1 XNOR_1_3_NUM24 (.ZN (XNOR_1_3_NUM24_OUT), .A1 (XNOR_1_1_NUM24_OUT), .A2 (XNOR_1_2_NUM24_OUT));
       NOR2_X1 XNOR_1_4_NUM24 (.ZN (N165), .A1 (XNOR_1_3_NUM24_OUT), .A2 (GND));
       wire XNOR_1_1_NUM25_OUT, XNOR_1_2_NUM25_OUT, XNOR_1_3_NUM25_OUT;
       NOR2_X1 XNOR_1_1_NUM25 (.ZN (XNOR_1_1_NUM25_OUT), .A1 (N134), .A2 (GND));
       NOR2_X1 XNOR_1_2_NUM25 (.ZN (XNOR_1_2_NUM25_OUT), .A1 (GND), .A2 (N56));
       NOR2_X1 XNOR_1_3_NUM25 (.ZN (XNOR_1_3_NUM25_OUT), .A1 (XNOR_1_1_NUM25_OUT), .A2 (XNOR_1_2_NUM25_OUT));
       NOR2_X1 XNOR_1_4_NUM25 (.ZN (N168), .A1 (XNOR_1_3_NUM25_OUT), .A2 (GND));
       wire XNOR_1_1_NUM26_OUT, XNOR_1_2_NUM26_OUT, XNOR_1_3_NUM26_OUT;
       NOR2_X1 XNOR_1_1_NUM26 (.ZN (XNOR_1_1_NUM26_OUT), .A1 (N138), .A2 (GND));
       NOR2_X1 XNOR_1_2_NUM26 (.ZN (XNOR_1_2_NUM26_OUT), .A1 (GND), .A2 (N69));
       NOR2_X1 XNOR_1_3_NUM26 (.ZN (XNOR_1_3_NUM26_OUT), .A1 (XNOR_1_1_NUM26_OUT), .A2 (XNOR_1_2_NUM26_OUT));
       NOR2_X1 XNOR_1_4_NUM26 (.ZN (N171), .A1 (XNOR_1_3_NUM26_OUT), .A2 (GND));
       wire XNOR_1_1_NUM27_OUT, XNOR_1_2_NUM27_OUT, XNOR_1_3_NUM27_OUT;
       NOR2_X1 XNOR_1_1_NUM27 (.ZN (XNOR_1_1_NUM27_OUT), .A1 (N142), .A2 (GND));
       NOR2_X1 XNOR_1_2_NUM27 (.ZN (XNOR_1_2_NUM27_OUT), .A1 (GND), .A2 (N82));
       NOR2_X1 XNOR_1_3_NUM27 (.ZN (XNOR_1_3_NUM27_OUT), .A1 (XNOR_1_1_NUM27_OUT), .A2 (XNOR_1_2_NUM27_OUT));
       NOR2_X1 XNOR_1_4_NUM27 (.ZN (N174), .A1 (XNOR_1_3_NUM27_OUT), .A2 (GND));
       wire XNOR_1_1_NUM28_OUT, XNOR_1_2_NUM28_OUT, XNOR_1_3_NUM28_OUT;
       NOR2_X1 XNOR_1_1_NUM28 (.ZN (XNOR_1_1_NUM28_OUT), .A1 (N146), .A2 (GND));
       NOR2_X1 XNOR_1_2_NUM28 (.ZN (XNOR_1_2_NUM28_OUT), .A1 (GND), .A2 (N95));
       NOR2_X1 XNOR_1_3_NUM28 (.ZN (XNOR_1_3_NUM28_OUT), .A1 (XNOR_1_1_NUM28_OUT), .A2 (XNOR_1_2_NUM28_OUT));
       NOR2_X1 XNOR_1_4_NUM28 (.ZN (N177), .A1 (XNOR_1_3_NUM28_OUT), .A2 (GND));
       wire XNOR_1_1_NUM29_OUT, XNOR_1_2_NUM29_OUT, XNOR_1_3_NUM29_OUT;
       NOR2_X1 XNOR_1_1_NUM29 (.ZN (XNOR_1_1_NUM29_OUT), .A1 (N150), .A2 (GND));
       NOR2_X1 XNOR_1_2_NUM29 (.ZN (XNOR_1_2_NUM29_OUT), .A1 (GND), .A2 (N108));
       NOR2_X1 XNOR_1_3_NUM29 (.ZN (XNOR_1_3_NUM29_OUT), .A1 (XNOR_1_1_NUM29_OUT), .A2 (XNOR_1_2_NUM29_OUT));
       NOR2_X1 XNOR_1_4_NUM29 (.ZN (N180), .A1 (XNOR_1_3_NUM29_OUT), .A2 (GND));
       NOR2_X1 XNOR_NUM30 (.ZN (N183), .A1 (N21), .A2 (N123));
       NOR2_X1 XNOR_NUM31 (.ZN (N184), .A1 (N27), .A2 (N123));
       NOR2_X1 XNOR_NUM32 (.ZN (N185), .A1 (N34), .A2 (N127));
       NOR2_X1 XNOR_NUM33 (.ZN (N186), .A1 (N40), .A2 (N127));
       NOR2_X1 XNOR_NUM34 (.ZN (N187), .A1 (N47), .A2 (N131));
       NOR2_X1 XNOR_NUM35 (.ZN (N188), .A1 (N53), .A2 (N131));
       NOR2_X1 XNOR_NUM36 (.ZN (N189), .A1 (N60), .A2 (N135));
       NOR2_X1 XNOR_NUM37 (.ZN (N190), .A1 (N66), .A2 (N135));
       NOR2_X1 XNOR_NUM38 (.ZN (N191), .A1 (N73), .A2 (N139));
       NOR2_X1 XNOR_NUM39 (.ZN (N192), .A1 (N79), .A2 (N139));
       NOR2_X1 XNOR_NUM40 (.ZN (N193), .A1 (N86), .A2 (N143));
       NOR2_X1 XNOR_NUM41 (.ZN (N194), .A1 (N92), .A2 (N143));
       NOR2_X1 XNOR_NUM42 (.ZN (N195), .A1 (N99), .A2 (N147));
       NOR2_X1 XNOR_NUM43 (.ZN (N196), .A1 (N105), .A2 (N147));
       NOR2_X1 XNOR_NUM44 (.ZN (N197), .A1 (N112), .A2 (N151));
       NOR2_X1 XNOR_NUM45 (.ZN (N198), .A1 (N115), .A2 (N151));
       wire XNOR_1_1_NUM46_OUT, XNOR_1_2_NUM46_OUT, XNOR_1_3_NUM46_OUT;
       NOR2_X1 XNOR_1_1_NUM46 (.ZN (XNOR_1_1_NUM46_OUT), .A1 (N154), .A2 (GND));
       NOR2_X1 XNOR_1_2_NUM46 (.ZN (XNOR_1_2_NUM46_OUT), .A1 (GND), .A2 (N159));
       NOR2_X1 XNOR_1_3_NUM46 (.ZN (XNOR_1_3_NUM46_OUT), .A1 (XNOR_1_1_NUM46_OUT), .A2 (XNOR_1_2_NUM46_OUT));

       wire XNOR_2_1_NUM46_OUT, XNOR_2_2_NUM46_OUT, XNOR_2_3_NUM46_OUT;
       NOR2_X1 XNOR_2_1_NUM46 (.ZN (XNOR_2_1_NUM46_OUT), .A1 (N162), .A2 (GND));
       NOR2_X1 XNOR_2_2_NUM46 (.ZN (XNOR_2_2_NUM46_OUT), .A1 (GND), .A2 (N165));
       NOR2_X1 XNOR_2_3_NUM46 (.ZN (XNOR_2_3_NUM46_OUT), .A1 (XNOR_2_1_NUM46_OUT), .A2 (XNOR_2_2_NUM46_OUT));

       wire XNOR_3_1_NUM46_OUT, XNOR_3_2_NUM46_OUT, XNOR_3_3_NUM46_OUT;
       NOR2_X1 XNOR_3_1_NUM46 (.ZN (XNOR_3_1_NUM46_OUT), .A1 (N168), .A2 (GND));
       NOR2_X1 XNOR_3_2_NUM46 (.ZN (XNOR_3_2_NUM46_OUT), .A1 (GND), .A2 (N171));
       NOR2_X1 XNOR_3_3_NUM46 (.ZN (XNOR_3_3_NUM46_OUT), .A1 (XNOR_3_1_NUM46_OUT), .A2 (XNOR_3_2_NUM46_OUT));

       wire XNOR_4_1_NUM46_OUT, XNOR_4_2_NUM46_OUT, XNOR_4_3_NUM46_OUT;
       NOR2_X1 XNOR_4_1_NUM46 (.ZN (XNOR_4_1_NUM46_OUT), .A1 (N174), .A2 (GND));
       NOR2_X1 XNOR_4_2_NUM46 (.ZN (XNOR_4_2_NUM46_OUT), .A1 (GND), .A2 (N177));
       NOR2_X1 XNOR_4_3_NUM46 (.ZN (XNOR_4_3_NUM46_OUT), .A1 (XNOR_4_1_NUM46_OUT), .A2 (XNOR_4_2_NUM46_OUT));

       wire XNOR_5_1_NUM46_OUT, XNOR_5_2_NUM46_OUT, XNOR_5_3_NUM46_OUT;
       NOR2_X1 XNOR_5_1_NUM46 (.ZN (XNOR_5_1_NUM46_OUT), .A1 (XNOR_1_3_NUM46_OUT), .A2 (GND));
       NOR2_X1 XNOR_5_2_NUM46 (.ZN (XNOR_5_2_NUM46_OUT), .A1 (GND), .A2 (XNOR_2_3_NUM46_OUT));
       NOR2_X1 XNOR_5_3_NUM46 (.ZN (XNOR_5_3_NUM46_OUT), .A1 (XNOR_5_1_NUM46_OUT), .A2 (XNOR_5_2_NUM46_OUT));

       wire XNOR_6_1_NUM46_OUT, XNOR_6_2_NUM46_OUT, XNOR_6_3_NUM46_OUT;
       NOR2_X1 XNOR_6_1_NUM46 (.ZN (XNOR_6_1_NUM46_OUT), .A1 (XNOR_3_3_NUM46_OUT), .A2 (GND));
       NOR2_X1 XNOR_6_2_NUM46 (.ZN (XNOR_6_2_NUM46_OUT), .A1 (GND), .A2 (XNOR_4_3_NUM46_OUT));
       NOR2_X1 XNOR_6_3_NUM46 (.ZN (XNOR_6_3_NUM46_OUT), .A1 (XNOR_6_1_NUM46_OUT), .A2 (XNOR_6_2_NUM46_OUT));

       wire XNOR_7_1_NUM46_OUT, XNOR_7_2_NUM46_OUT, XNOR_7_3_NUM46_OUT;
       NOR2_X1 XNOR_7_1_NUM46 (.ZN (XNOR_7_1_NUM46_OUT), .A1 (XNOR_5_3_NUM46_OUT), .A2 (GND));
       NOR2_X1 XNOR_7_2_NUM46 (.ZN (XNOR_7_2_NUM46_OUT), .A1 (GND), .A2 (XNOR_6_3_NUM46_OUT));
       NOR2_X1 XNOR_7_3_NUM46 (.ZN (XNOR_7_3_NUM46_OUT), .A1 (XNOR_7_1_NUM46_OUT), .A2 (XNOR_7_2_NUM46_OUT));

       wire XNOR_8_1_NUM46_OUT, XNOR_8_2_NUM46_OUT, XNOR_8_3_NUM46_OUT;
       NOR2_X1 XNOR_8_1_NUM46 (.ZN (XNOR_8_1_NUM46_OUT), .A1 (XNOR_7_3_NUM46_OUT), .A2 (GND));
       NOR2_X1 XNOR_8_2_NUM46 (.ZN (XNOR_8_2_NUM46_OUT), .A1 (GND), .A2 (N180));
       NOR2_X1 XNOR_8_3_NUM46 (.ZN (N199), .A1 (XNOR_8_1_NUM46_OUT), .A2 (XNOR_8_2_NUM46_OUT));
       NOR2_X1 XNOR_NUM47 (.ZN (N203), .A1 (N199), .A2 (GND));
       NOR2_X1 XNOR_NUM48 (.ZN (N213), .A1 (N199), .A2 (GND));
       NOR2_X1 XNOR_NUM49 (.ZN (N223), .A1 (N199), .A2 (GND));
       wire XNOR_1_1_NUM50_OUT, XNOR_1_2_NUM50_OUT, XNOR_1_3_NUM50_OUT, XNOR_1_4_NUM50_OUT;
       NOR2_X1 XNOR_1_1_NUM50 (.ZN (XNOR_1_1_NUM50_OUT), .A1 (N203), .A2 (GND));
       NOR2_X1 XNOR_1_2_NUM50 (.ZN (XNOR_1_2_NUM50_OUT), .A1 (GND), .A2 (N154));
       NOR2_X1 XNOR_1_3_NUM50 (.ZN (XNOR_1_3_NUM50_OUT), .A1 (XNOR_1_1_NUM50_OUT), .A2 (XNOR_1_2_NUM50_OUT));
       NOR2_X1 XNOR_1_4_NUM50 (.ZN (XNOR_1_4_NUM50_OUT), .A1 (N203), .A2 (N154));
       NOR2_X1 XNOR_1_5_NUM50 (.ZN (N224), .A1 (XNOR_1_3_NUM50_OUT), .A2 (XNOR_1_4_NUM50_OUT));
       wire XNOR_1_1_NUM51_OUT, XNOR_1_2_NUM51_OUT, XNOR_1_3_NUM51_OUT, XNOR_1_4_NUM51_OUT;
       NOR2_X1 XNOR_1_1_NUM51 (.ZN (XNOR_1_1_NUM51_OUT), .A1 (N203), .A2 (GND));
       NOR2_X1 XNOR_1_2_NUM51 (.ZN (XNOR_1_2_NUM51_OUT), .A1 (GND), .A2 (N159));
       NOR2_X1 XNOR_1_3_NUM51 (.ZN (XNOR_1_3_NUM51_OUT), .A1 (XNOR_1_1_NUM51_OUT), .A2 (XNOR_1_2_NUM51_OUT));
       NOR2_X1 XNOR_1_4_NUM51 (.ZN (XNOR_1_4_NUM51_OUT), .A1 (N203), .A2 (N159));
       NOR2_X1 XNOR_1_5_NUM51 (.ZN (N227), .A1 (XNOR_1_3_NUM51_OUT), .A2 (XNOR_1_4_NUM51_OUT));
       wire XNOR_1_1_NUM52_OUT, XNOR_1_2_NUM52_OUT, XNOR_1_3_NUM52_OUT, XNOR_1_4_NUM52_OUT;
       NOR2_X1 XNOR_1_1_NUM52 (.ZN (XNOR_1_1_NUM52_OUT), .A1 (N203), .A2 (GND));
       NOR2_X1 XNOR_1_2_NUM52 (.ZN (XNOR_1_2_NUM52_OUT), .A1 (GND), .A2 (N162));
       NOR2_X1 XNOR_1_3_NUM52 (.ZN (XNOR_1_3_NUM52_OUT), .A1 (XNOR_1_1_NUM52_OUT), .A2 (XNOR_1_2_NUM52_OUT));
       NOR2_X1 XNOR_1_4_NUM52 (.ZN (XNOR_1_4_NUM52_OUT), .A1 (N203), .A2 (N162));
       NOR2_X1 XNOR_1_5_NUM52 (.ZN (N230), .A1 (XNOR_1_3_NUM52_OUT), .A2 (XNOR_1_4_NUM52_OUT));
       wire XNOR_1_1_NUM53_OUT, XNOR_1_2_NUM53_OUT, XNOR_1_3_NUM53_OUT, XNOR_1_4_NUM53_OUT;
       NOR2_X1 XNOR_1_1_NUM53 (.ZN (XNOR_1_1_NUM53_OUT), .A1 (N203), .A2 (GND));
       NOR2_X1 XNOR_1_2_NUM53 (.ZN (XNOR_1_2_NUM53_OUT), .A1 (GND), .A2 (N165));
       NOR2_X1 XNOR_1_3_NUM53 (.ZN (XNOR_1_3_NUM53_OUT), .A1 (XNOR_1_1_NUM53_OUT), .A2 (XNOR_1_2_NUM53_OUT));
       NOR2_X1 XNOR_1_4_NUM53 (.ZN (XNOR_1_4_NUM53_OUT), .A1 (N203), .A2 (N165));
       NOR2_X1 XNOR_1_5_NUM53 (.ZN (N233), .A1 (XNOR_1_3_NUM53_OUT), .A2 (XNOR_1_4_NUM53_OUT));
       wire XNOR_1_1_NUM54_OUT, XNOR_1_2_NUM54_OUT, XNOR_1_3_NUM54_OUT, XNOR_1_4_NUM54_OUT;
       NOR2_X1 XNOR_1_1_NUM54 (.ZN (XNOR_1_1_NUM54_OUT), .A1 (N203), .A2 (GND));
       NOR2_X1 XNOR_1_2_NUM54 (.ZN (XNOR_1_2_NUM54_OUT), .A1 (GND), .A2 (N168));
       NOR2_X1 XNOR_1_3_NUM54 (.ZN (XNOR_1_3_NUM54_OUT), .A1 (XNOR_1_1_NUM54_OUT), .A2 (XNOR_1_2_NUM54_OUT));
       NOR2_X1 XNOR_1_4_NUM54 (.ZN (XNOR_1_4_NUM54_OUT), .A1 (N203), .A2 (N168));
       NOR2_X1 XNOR_1_5_NUM54 (.ZN (N236), .A1 (XNOR_1_3_NUM54_OUT), .A2 (XNOR_1_4_NUM54_OUT));
       wire XNOR_1_1_NUM55_OUT, XNOR_1_2_NUM55_OUT, XNOR_1_3_NUM55_OUT, XNOR_1_4_NUM55_OUT;
       NOR2_X1 XNOR_1_1_NUM55 (.ZN (XNOR_1_1_NUM55_OUT), .A1 (N203), .A2 (GND));
       NOR2_X1 XNOR_1_2_NUM55 (.ZN (XNOR_1_2_NUM55_OUT), .A1 (GND), .A2 (N171));
       NOR2_X1 XNOR_1_3_NUM55 (.ZN (XNOR_1_3_NUM55_OUT), .A1 (XNOR_1_1_NUM55_OUT), .A2 (XNOR_1_2_NUM55_OUT));
       NOR2_X1 XNOR_1_4_NUM55 (.ZN (XNOR_1_4_NUM55_OUT), .A1 (N203), .A2 (N171));
       NOR2_X1 XNOR_1_5_NUM55 (.ZN (N239), .A1 (XNOR_1_3_NUM55_OUT), .A2 (XNOR_1_4_NUM55_OUT));
       wire XNOR_1_1_NUM56_OUT, XNOR_1_2_NUM56_OUT, XNOR_1_3_NUM56_OUT;
       NOR2_X1 XNOR_1_1_NUM56 (.ZN (XNOR_1_1_NUM56_OUT), .A1 (N1), .A2 (GND));
       NOR2_X1 XNOR_1_2_NUM56 (.ZN (XNOR_1_2_NUM56_OUT), .A1 (GND), .A2 (N213));
       NOR2_X1 XNOR_1_3_NUM56 (.ZN (XNOR_1_3_NUM56_OUT), .A1 (XNOR_1_1_NUM56_OUT), .A2 (XNOR_1_2_NUM56_OUT));
       NOR2_X1 XNOR_1_4_NUM56 (.ZN (N242), .A1 (XNOR_1_3_NUM56_OUT), .A2 (GND));
       wire XNOR_1_1_NUM57_OUT, XNOR_1_2_NUM57_OUT, XNOR_1_3_NUM57_OUT, XNOR_1_4_NUM57_OUT;
       NOR2_X1 XNOR_1_1_NUM57 (.ZN (XNOR_1_1_NUM57_OUT), .A1 (N203), .A2 (GND));
       NOR2_X1 XNOR_1_2_NUM57 (.ZN (XNOR_1_2_NUM57_OUT), .A1 (GND), .A2 (N174));
       NOR2_X1 XNOR_1_3_NUM57 (.ZN (XNOR_1_3_NUM57_OUT), .A1 (XNOR_1_1_NUM57_OUT), .A2 (XNOR_1_2_NUM57_OUT));
       NOR2_X1 XNOR_1_4_NUM57 (.ZN (XNOR_1_4_NUM57_OUT), .A1 (N203), .A2 (N174));
       NOR2_X1 XNOR_1_5_NUM57 (.ZN (N243), .A1 (XNOR_1_3_NUM57_OUT), .A2 (XNOR_1_4_NUM57_OUT));
       wire XNOR_1_1_NUM58_OUT, XNOR_1_2_NUM58_OUT, XNOR_1_3_NUM58_OUT;
       NOR2_X1 XNOR_1_1_NUM58 (.ZN (XNOR_1_1_NUM58_OUT), .A1 (N213), .A2 (GND));
       NOR2_X1 XNOR_1_2_NUM58 (.ZN (XNOR_1_2_NUM58_OUT), .A1 (GND), .A2 (N11));
       NOR2_X1 XNOR_1_3_NUM58 (.ZN (XNOR_1_3_NUM58_OUT), .A1 (XNOR_1_1_NUM58_OUT), .A2 (XNOR_1_2_NUM58_OUT));
       NOR2_X1 XNOR_1_4_NUM58 (.ZN (N246), .A1 (XNOR_1_3_NUM58_OUT), .A2 (GND));
       wire XNOR_1_1_NUM59_OUT, XNOR_1_2_NUM59_OUT, XNOR_1_3_NUM59_OUT, XNOR_1_4_NUM59_OUT;
       NOR2_X1 XNOR_1_1_NUM59 (.ZN (XNOR_1_1_NUM59_OUT), .A1 (N203), .A2 (GND));
       NOR2_X1 XNOR_1_2_NUM59 (.ZN (XNOR_1_2_NUM59_OUT), .A1 (GND), .A2 (N177));
       NOR2_X1 XNOR_1_3_NUM59 (.ZN (XNOR_1_3_NUM59_OUT), .A1 (XNOR_1_1_NUM59_OUT), .A2 (XNOR_1_2_NUM59_OUT));
       NOR2_X1 XNOR_1_4_NUM59 (.ZN (XNOR_1_4_NUM59_OUT), .A1 (N203), .A2 (N177));
       NOR2_X1 XNOR_1_5_NUM59 (.ZN (N247), .A1 (XNOR_1_3_NUM59_OUT), .A2 (XNOR_1_4_NUM59_OUT));
       wire XNOR_1_1_NUM60_OUT, XNOR_1_2_NUM60_OUT, XNOR_1_3_NUM60_OUT;
       NOR2_X1 XNOR_1_1_NUM60 (.ZN (XNOR_1_1_NUM60_OUT), .A1 (N213), .A2 (GND));
       NOR2_X1 XNOR_1_2_NUM60 (.ZN (XNOR_1_2_NUM60_OUT), .A1 (GND), .A2 (N24));
       NOR2_X1 XNOR_1_3_NUM60 (.ZN (XNOR_1_3_NUM60_OUT), .A1 (XNOR_1_1_NUM60_OUT), .A2 (XNOR_1_2_NUM60_OUT));
       NOR2_X1 XNOR_1_4_NUM60 (.ZN (N250), .A1 (XNOR_1_3_NUM60_OUT), .A2 (GND));
       wire XNOR_1_1_NUM61_OUT, XNOR_1_2_NUM61_OUT, XNOR_1_3_NUM61_OUT, XNOR_1_4_NUM61_OUT;
       NOR2_X1 XNOR_1_1_NUM61 (.ZN (XNOR_1_1_NUM61_OUT), .A1 (N203), .A2 (GND));
       NOR2_X1 XNOR_1_2_NUM61 (.ZN (XNOR_1_2_NUM61_OUT), .A1 (GND), .A2 (N180));
       NOR2_X1 XNOR_1_3_NUM61 (.ZN (XNOR_1_3_NUM61_OUT), .A1 (XNOR_1_1_NUM61_OUT), .A2 (XNOR_1_2_NUM61_OUT));
       NOR2_X1 XNOR_1_4_NUM61 (.ZN (XNOR_1_4_NUM61_OUT), .A1 (N203), .A2 (N180));
       NOR2_X1 XNOR_1_5_NUM61 (.ZN (N251), .A1 (XNOR_1_3_NUM61_OUT), .A2 (XNOR_1_4_NUM61_OUT));
       wire XNOR_1_1_NUM62_OUT, XNOR_1_2_NUM62_OUT, XNOR_1_3_NUM62_OUT;
       NOR2_X1 XNOR_1_1_NUM62 (.ZN (XNOR_1_1_NUM62_OUT), .A1 (N213), .A2 (GND));
       NOR2_X1 XNOR_1_2_NUM62 (.ZN (XNOR_1_2_NUM62_OUT), .A1 (GND), .A2 (N37));
       NOR2_X1 XNOR_1_3_NUM62 (.ZN (XNOR_1_3_NUM62_OUT), .A1 (XNOR_1_1_NUM62_OUT), .A2 (XNOR_1_2_NUM62_OUT));
       NOR2_X1 XNOR_1_4_NUM62 (.ZN (N254), .A1 (XNOR_1_3_NUM62_OUT), .A2 (GND));
       wire XNOR_1_1_NUM63_OUT, XNOR_1_2_NUM63_OUT, XNOR_1_3_NUM63_OUT;
       NOR2_X1 XNOR_1_1_NUM63 (.ZN (XNOR_1_1_NUM63_OUT), .A1 (N213), .A2 (GND));
       NOR2_X1 XNOR_1_2_NUM63 (.ZN (XNOR_1_2_NUM63_OUT), .A1 (GND), .A2 (N50));
       NOR2_X1 XNOR_1_3_NUM63 (.ZN (XNOR_1_3_NUM63_OUT), .A1 (XNOR_1_1_NUM63_OUT), .A2 (XNOR_1_2_NUM63_OUT));
       NOR2_X1 XNOR_1_4_NUM63 (.ZN (N255), .A1 (XNOR_1_3_NUM63_OUT), .A2 (GND));
       wire XNOR_1_1_NUM64_OUT, XNOR_1_2_NUM64_OUT, XNOR_1_3_NUM64_OUT;
       NOR2_X1 XNOR_1_1_NUM64 (.ZN (XNOR_1_1_NUM64_OUT), .A1 (N213), .A2 (GND));
       NOR2_X1 XNOR_1_2_NUM64 (.ZN (XNOR_1_2_NUM64_OUT), .A1 (GND), .A2 (N63));
       NOR2_X1 XNOR_1_3_NUM64 (.ZN (XNOR_1_3_NUM64_OUT), .A1 (XNOR_1_1_NUM64_OUT), .A2 (XNOR_1_2_NUM64_OUT));
       NOR2_X1 XNOR_1_4_NUM64 (.ZN (N256), .A1 (XNOR_1_3_NUM64_OUT), .A2 (GND));
       wire XNOR_1_1_NUM65_OUT, XNOR_1_2_NUM65_OUT, XNOR_1_3_NUM65_OUT;
       NOR2_X1 XNOR_1_1_NUM65 (.ZN (XNOR_1_1_NUM65_OUT), .A1 (N213), .A2 (GND));
       NOR2_X1 XNOR_1_2_NUM65 (.ZN (XNOR_1_2_NUM65_OUT), .A1 (GND), .A2 (N76));
       NOR2_X1 XNOR_1_3_NUM65 (.ZN (XNOR_1_3_NUM65_OUT), .A1 (XNOR_1_1_NUM65_OUT), .A2 (XNOR_1_2_NUM65_OUT));
       NOR2_X1 XNOR_1_4_NUM65 (.ZN (N257), .A1 (XNOR_1_3_NUM65_OUT), .A2 (GND));
       wire XNOR_1_1_NUM66_OUT, XNOR_1_2_NUM66_OUT, XNOR_1_3_NUM66_OUT;
       NOR2_X1 XNOR_1_1_NUM66 (.ZN (XNOR_1_1_NUM66_OUT), .A1 (N213), .A2 (GND));
       NOR2_X1 XNOR_1_2_NUM66 (.ZN (XNOR_1_2_NUM66_OUT), .A1 (GND), .A2 (N89));
       NOR2_X1 XNOR_1_3_NUM66 (.ZN (XNOR_1_3_NUM66_OUT), .A1 (XNOR_1_1_NUM66_OUT), .A2 (XNOR_1_2_NUM66_OUT));
       NOR2_X1 XNOR_1_4_NUM66 (.ZN (N258), .A1 (XNOR_1_3_NUM66_OUT), .A2 (GND));
       wire XNOR_1_1_NUM67_OUT, XNOR_1_2_NUM67_OUT, XNOR_1_3_NUM67_OUT;
       NOR2_X1 XNOR_1_1_NUM67 (.ZN (XNOR_1_1_NUM67_OUT), .A1 (N213), .A2 (GND));
       NOR2_X1 XNOR_1_2_NUM67 (.ZN (XNOR_1_2_NUM67_OUT), .A1 (GND), .A2 (N102));
       NOR2_X1 XNOR_1_3_NUM67 (.ZN (XNOR_1_3_NUM67_OUT), .A1 (XNOR_1_1_NUM67_OUT), .A2 (XNOR_1_2_NUM67_OUT));
       NOR2_X1 XNOR_1_4_NUM67 (.ZN (N259), .A1 (XNOR_1_3_NUM67_OUT), .A2 (GND));
       wire XNOR_1_1_NUM68_OUT, XNOR_1_2_NUM68_OUT, XNOR_1_3_NUM68_OUT;
       NOR2_X1 XNOR_1_1_NUM68 (.ZN (XNOR_1_1_NUM68_OUT), .A1 (N224), .A2 (GND));
       NOR2_X1 XNOR_1_2_NUM68 (.ZN (XNOR_1_2_NUM68_OUT), .A1 (GND), .A2 (N157));
       NOR2_X1 XNOR_1_3_NUM68 (.ZN (XNOR_1_3_NUM68_OUT), .A1 (XNOR_1_1_NUM68_OUT), .A2 (XNOR_1_2_NUM68_OUT));
       NOR2_X1 XNOR_1_4_NUM68 (.ZN (N260), .A1 (XNOR_1_3_NUM68_OUT), .A2 (GND));
       wire XNOR_1_1_NUM69_OUT, XNOR_1_2_NUM69_OUT, XNOR_1_3_NUM69_OUT;
       NOR2_X1 XNOR_1_1_NUM69 (.ZN (XNOR_1_1_NUM69_OUT), .A1 (N224), .A2 (GND));
       NOR2_X1 XNOR_1_2_NUM69 (.ZN (XNOR_1_2_NUM69_OUT), .A1 (GND), .A2 (N158));
       NOR2_X1 XNOR_1_3_NUM69 (.ZN (XNOR_1_3_NUM69_OUT), .A1 (XNOR_1_1_NUM69_OUT), .A2 (XNOR_1_2_NUM69_OUT));
       NOR2_X1 XNOR_1_4_NUM69 (.ZN (N263), .A1 (XNOR_1_3_NUM69_OUT), .A2 (GND));
       wire XNOR_1_1_NUM70_OUT, XNOR_1_2_NUM70_OUT, XNOR_1_3_NUM70_OUT;
       NOR2_X1 XNOR_1_1_NUM70 (.ZN (XNOR_1_1_NUM70_OUT), .A1 (N227), .A2 (GND));
       NOR2_X1 XNOR_1_2_NUM70 (.ZN (XNOR_1_2_NUM70_OUT), .A1 (GND), .A2 (N183));
       NOR2_X1 XNOR_1_3_NUM70 (.ZN (XNOR_1_3_NUM70_OUT), .A1 (XNOR_1_1_NUM70_OUT), .A2 (XNOR_1_2_NUM70_OUT));
       NOR2_X1 XNOR_1_4_NUM70 (.ZN (N264), .A1 (XNOR_1_3_NUM70_OUT), .A2 (GND));
       wire XNOR_1_1_NUM71_OUT, XNOR_1_2_NUM71_OUT, XNOR_1_3_NUM71_OUT;
       NOR2_X1 XNOR_1_1_NUM71 (.ZN (XNOR_1_1_NUM71_OUT), .A1 (N230), .A2 (GND));
       NOR2_X1 XNOR_1_2_NUM71 (.ZN (XNOR_1_2_NUM71_OUT), .A1 (GND), .A2 (N185));
       NOR2_X1 XNOR_1_3_NUM71 (.ZN (XNOR_1_3_NUM71_OUT), .A1 (XNOR_1_1_NUM71_OUT), .A2 (XNOR_1_2_NUM71_OUT));
       NOR2_X1 XNOR_1_4_NUM71 (.ZN (N267), .A1 (XNOR_1_3_NUM71_OUT), .A2 (GND));
       wire XNOR_1_1_NUM72_OUT, XNOR_1_2_NUM72_OUT, XNOR_1_3_NUM72_OUT;
       NOR2_X1 XNOR_1_1_NUM72 (.ZN (XNOR_1_1_NUM72_OUT), .A1 (N233), .A2 (GND));
       NOR2_X1 XNOR_1_2_NUM72 (.ZN (XNOR_1_2_NUM72_OUT), .A1 (GND), .A2 (N187));
       NOR2_X1 XNOR_1_3_NUM72 (.ZN (XNOR_1_3_NUM72_OUT), .A1 (XNOR_1_1_NUM72_OUT), .A2 (XNOR_1_2_NUM72_OUT));
       NOR2_X1 XNOR_1_4_NUM72 (.ZN (N270), .A1 (XNOR_1_3_NUM72_OUT), .A2 (GND));
       wire XNOR_1_1_NUM73_OUT, XNOR_1_2_NUM73_OUT, XNOR_1_3_NUM73_OUT;
       NOR2_X1 XNOR_1_1_NUM73 (.ZN (XNOR_1_1_NUM73_OUT), .A1 (N236), .A2 (GND));
       NOR2_X1 XNOR_1_2_NUM73 (.ZN (XNOR_1_2_NUM73_OUT), .A1 (GND), .A2 (N189));
       NOR2_X1 XNOR_1_3_NUM73 (.ZN (XNOR_1_3_NUM73_OUT), .A1 (XNOR_1_1_NUM73_OUT), .A2 (XNOR_1_2_NUM73_OUT));
       NOR2_X1 XNOR_1_4_NUM73 (.ZN (N273), .A1 (XNOR_1_3_NUM73_OUT), .A2 (GND));
       wire XNOR_1_1_NUM74_OUT, XNOR_1_2_NUM74_OUT, XNOR_1_3_NUM74_OUT;
       NOR2_X1 XNOR_1_1_NUM74 (.ZN (XNOR_1_1_NUM74_OUT), .A1 (N239), .A2 (GND));
       NOR2_X1 XNOR_1_2_NUM74 (.ZN (XNOR_1_2_NUM74_OUT), .A1 (GND), .A2 (N191));
       NOR2_X1 XNOR_1_3_NUM74 (.ZN (XNOR_1_3_NUM74_OUT), .A1 (XNOR_1_1_NUM74_OUT), .A2 (XNOR_1_2_NUM74_OUT));
       NOR2_X1 XNOR_1_4_NUM74 (.ZN (N276), .A1 (XNOR_1_3_NUM74_OUT), .A2 (GND));
       wire XNOR_1_1_NUM75_OUT, XNOR_1_2_NUM75_OUT, XNOR_1_3_NUM75_OUT;
       NOR2_X1 XNOR_1_1_NUM75 (.ZN (XNOR_1_1_NUM75_OUT), .A1 (N243), .A2 (GND));
       NOR2_X1 XNOR_1_2_NUM75 (.ZN (XNOR_1_2_NUM75_OUT), .A1 (GND), .A2 (N193));
       NOR2_X1 XNOR_1_3_NUM75 (.ZN (XNOR_1_3_NUM75_OUT), .A1 (XNOR_1_1_NUM75_OUT), .A2 (XNOR_1_2_NUM75_OUT));
       NOR2_X1 XNOR_1_4_NUM75 (.ZN (N279), .A1 (XNOR_1_3_NUM75_OUT), .A2 (GND));
       wire XNOR_1_1_NUM76_OUT, XNOR_1_2_NUM76_OUT, XNOR_1_3_NUM76_OUT;
       NOR2_X1 XNOR_1_1_NUM76 (.ZN (XNOR_1_1_NUM76_OUT), .A1 (N247), .A2 (GND));
       NOR2_X1 XNOR_1_2_NUM76 (.ZN (XNOR_1_2_NUM76_OUT), .A1 (GND), .A2 (N195));
       NOR2_X1 XNOR_1_3_NUM76 (.ZN (XNOR_1_3_NUM76_OUT), .A1 (XNOR_1_1_NUM76_OUT), .A2 (XNOR_1_2_NUM76_OUT));
       NOR2_X1 XNOR_1_4_NUM76 (.ZN (N282), .A1 (XNOR_1_3_NUM76_OUT), .A2 (GND));
       wire XNOR_1_1_NUM77_OUT, XNOR_1_2_NUM77_OUT, XNOR_1_3_NUM77_OUT;
       NOR2_X1 XNOR_1_1_NUM77 (.ZN (XNOR_1_1_NUM77_OUT), .A1 (N251), .A2 (GND));
       NOR2_X1 XNOR_1_2_NUM77 (.ZN (XNOR_1_2_NUM77_OUT), .A1 (GND), .A2 (N197));
       NOR2_X1 XNOR_1_3_NUM77 (.ZN (XNOR_1_3_NUM77_OUT), .A1 (XNOR_1_1_NUM77_OUT), .A2 (XNOR_1_2_NUM77_OUT));
       NOR2_X1 XNOR_1_4_NUM77 (.ZN (N285), .A1 (XNOR_1_3_NUM77_OUT), .A2 (GND));
       wire XNOR_1_1_NUM78_OUT, XNOR_1_2_NUM78_OUT, XNOR_1_3_NUM78_OUT;
       NOR2_X1 XNOR_1_1_NUM78 (.ZN (XNOR_1_1_NUM78_OUT), .A1 (N227), .A2 (GND));
       NOR2_X1 XNOR_1_2_NUM78 (.ZN (XNOR_1_2_NUM78_OUT), .A1 (GND), .A2 (N184));
       NOR2_X1 XNOR_1_3_NUM78 (.ZN (XNOR_1_3_NUM78_OUT), .A1 (XNOR_1_1_NUM78_OUT), .A2 (XNOR_1_2_NUM78_OUT));
       NOR2_X1 XNOR_1_4_NUM78 (.ZN (N288), .A1 (XNOR_1_3_NUM78_OUT), .A2 (GND));
       wire XNOR_1_1_NUM79_OUT, XNOR_1_2_NUM79_OUT, XNOR_1_3_NUM79_OUT;
       NOR2_X1 XNOR_1_1_NUM79 (.ZN (XNOR_1_1_NUM79_OUT), .A1 (N230), .A2 (GND));
       NOR2_X1 XNOR_1_2_NUM79 (.ZN (XNOR_1_2_NUM79_OUT), .A1 (GND), .A2 (N186));
       NOR2_X1 XNOR_1_3_NUM79 (.ZN (XNOR_1_3_NUM79_OUT), .A1 (XNOR_1_1_NUM79_OUT), .A2 (XNOR_1_2_NUM79_OUT));
       NOR2_X1 XNOR_1_4_NUM79 (.ZN (N289), .A1 (XNOR_1_3_NUM79_OUT), .A2 (GND));
       wire XNOR_1_1_NUM80_OUT, XNOR_1_2_NUM80_OUT, XNOR_1_3_NUM80_OUT;
       NOR2_X1 XNOR_1_1_NUM80 (.ZN (XNOR_1_1_NUM80_OUT), .A1 (N233), .A2 (GND));
       NOR2_X1 XNOR_1_2_NUM80 (.ZN (XNOR_1_2_NUM80_OUT), .A1 (GND), .A2 (N188));
       NOR2_X1 XNOR_1_3_NUM80 (.ZN (XNOR_1_3_NUM80_OUT), .A1 (XNOR_1_1_NUM80_OUT), .A2 (XNOR_1_2_NUM80_OUT));
       NOR2_X1 XNOR_1_4_NUM80 (.ZN (N290), .A1 (XNOR_1_3_NUM80_OUT), .A2 (GND));
       wire XNOR_1_1_NUM81_OUT, XNOR_1_2_NUM81_OUT, XNOR_1_3_NUM81_OUT;
       NOR2_X1 XNOR_1_1_NUM81 (.ZN (XNOR_1_1_NUM81_OUT), .A1 (N236), .A2 (GND));
       NOR2_X1 XNOR_1_2_NUM81 (.ZN (XNOR_1_2_NUM81_OUT), .A1 (GND), .A2 (N190));
       NOR2_X1 XNOR_1_3_NUM81 (.ZN (XNOR_1_3_NUM81_OUT), .A1 (XNOR_1_1_NUM81_OUT), .A2 (XNOR_1_2_NUM81_OUT));
       NOR2_X1 XNOR_1_4_NUM81 (.ZN (N291), .A1 (XNOR_1_3_NUM81_OUT), .A2 (GND));
       wire XNOR_1_1_NUM82_OUT, XNOR_1_2_NUM82_OUT, XNOR_1_3_NUM82_OUT;
       NOR2_X1 XNOR_1_1_NUM82 (.ZN (XNOR_1_1_NUM82_OUT), .A1 (N239), .A2 (GND));
       NOR2_X1 XNOR_1_2_NUM82 (.ZN (XNOR_1_2_NUM82_OUT), .A1 (GND), .A2 (N192));
       NOR2_X1 XNOR_1_3_NUM82 (.ZN (XNOR_1_3_NUM82_OUT), .A1 (XNOR_1_1_NUM82_OUT), .A2 (XNOR_1_2_NUM82_OUT));
       NOR2_X1 XNOR_1_4_NUM82 (.ZN (N292), .A1 (XNOR_1_3_NUM82_OUT), .A2 (GND));
       wire XNOR_1_1_NUM83_OUT, XNOR_1_2_NUM83_OUT, XNOR_1_3_NUM83_OUT;
       NOR2_X1 XNOR_1_1_NUM83 (.ZN (XNOR_1_1_NUM83_OUT), .A1 (N243), .A2 (GND));
       NOR2_X1 XNOR_1_2_NUM83 (.ZN (XNOR_1_2_NUM83_OUT), .A1 (GND), .A2 (N194));
       NOR2_X1 XNOR_1_3_NUM83 (.ZN (XNOR_1_3_NUM83_OUT), .A1 (XNOR_1_1_NUM83_OUT), .A2 (XNOR_1_2_NUM83_OUT));
       NOR2_X1 XNOR_1_4_NUM83 (.ZN (N293), .A1 (XNOR_1_3_NUM83_OUT), .A2 (GND));
       wire XNOR_1_1_NUM84_OUT, XNOR_1_2_NUM84_OUT, XNOR_1_3_NUM84_OUT;
       NOR2_X1 XNOR_1_1_NUM84 (.ZN (XNOR_1_1_NUM84_OUT), .A1 (N247), .A2 (GND));
       NOR2_X1 XNOR_1_2_NUM84 (.ZN (XNOR_1_2_NUM84_OUT), .A1 (GND), .A2 (N196));
       NOR2_X1 XNOR_1_3_NUM84 (.ZN (XNOR_1_3_NUM84_OUT), .A1 (XNOR_1_1_NUM84_OUT), .A2 (XNOR_1_2_NUM84_OUT));
       NOR2_X1 XNOR_1_4_NUM84 (.ZN (N294), .A1 (XNOR_1_3_NUM84_OUT), .A2 (GND));
       wire XNOR_1_1_NUM85_OUT, XNOR_1_2_NUM85_OUT, XNOR_1_3_NUM85_OUT;
       NOR2_X1 XNOR_1_1_NUM85 (.ZN (XNOR_1_1_NUM85_OUT), .A1 (N251), .A2 (GND));
       NOR2_X1 XNOR_1_2_NUM85 (.ZN (XNOR_1_2_NUM85_OUT), .A1 (GND), .A2 (N198));
       NOR2_X1 XNOR_1_3_NUM85 (.ZN (XNOR_1_3_NUM85_OUT), .A1 (XNOR_1_1_NUM85_OUT), .A2 (XNOR_1_2_NUM85_OUT));
       NOR2_X1 XNOR_1_4_NUM85 (.ZN (N295), .A1 (XNOR_1_3_NUM85_OUT), .A2 (GND));
       wire XNOR_1_1_NUM86_OUT, XNOR_1_2_NUM86_OUT, XNOR_1_3_NUM86_OUT;
       NOR2_X1 XNOR_1_1_NUM86 (.ZN (XNOR_1_1_NUM86_OUT), .A1 (N260), .A2 (GND));
       NOR2_X1 XNOR_1_2_NUM86 (.ZN (XNOR_1_2_NUM86_OUT), .A1 (GND), .A2 (N264));
       NOR2_X1 XNOR_1_3_NUM86 (.ZN (XNOR_1_3_NUM86_OUT), .A1 (XNOR_1_1_NUM86_OUT), .A2 (XNOR_1_2_NUM86_OUT));

       wire XNOR_2_1_NUM86_OUT, XNOR_2_2_NUM86_OUT, XNOR_2_3_NUM86_OUT;
       NOR2_X1 XNOR_2_1_NUM86 (.ZN (XNOR_2_1_NUM86_OUT), .A1 (N267), .A2 (GND));
       NOR2_X1 XNOR_2_2_NUM86 (.ZN (XNOR_2_2_NUM86_OUT), .A1 (GND), .A2 (N270));
       NOR2_X1 XNOR_2_3_NUM86 (.ZN (XNOR_2_3_NUM86_OUT), .A1 (XNOR_2_1_NUM86_OUT), .A2 (XNOR_2_2_NUM86_OUT));

       wire XNOR_3_1_NUM86_OUT, XNOR_3_2_NUM86_OUT, XNOR_3_3_NUM86_OUT;
       NOR2_X1 XNOR_3_1_NUM86 (.ZN (XNOR_3_1_NUM86_OUT), .A1 (N273), .A2 (GND));
       NOR2_X1 XNOR_3_2_NUM86 (.ZN (XNOR_3_2_NUM86_OUT), .A1 (GND), .A2 (N276));
       NOR2_X1 XNOR_3_3_NUM86 (.ZN (XNOR_3_3_NUM86_OUT), .A1 (XNOR_3_1_NUM86_OUT), .A2 (XNOR_3_2_NUM86_OUT));

       wire XNOR_4_1_NUM86_OUT, XNOR_4_2_NUM86_OUT, XNOR_4_3_NUM86_OUT;
       NOR2_X1 XNOR_4_1_NUM86 (.ZN (XNOR_4_1_NUM86_OUT), .A1 (N279), .A2 (GND));
       NOR2_X1 XNOR_4_2_NUM86 (.ZN (XNOR_4_2_NUM86_OUT), .A1 (GND), .A2 (N282));
       NOR2_X1 XNOR_4_3_NUM86 (.ZN (XNOR_4_3_NUM86_OUT), .A1 (XNOR_4_1_NUM86_OUT), .A2 (XNOR_4_2_NUM86_OUT));

       wire XNOR_5_1_NUM86_OUT, XNOR_5_2_NUM86_OUT, XNOR_5_3_NUM86_OUT;
       NOR2_X1 XNOR_5_1_NUM86 (.ZN (XNOR_5_1_NUM86_OUT), .A1 (XNOR_1_3_NUM86_OUT), .A2 (GND));
       NOR2_X1 XNOR_5_2_NUM86 (.ZN (XNOR_5_2_NUM86_OUT), .A1 (GND), .A2 (XNOR_2_3_NUM86_OUT));
       NOR2_X1 XNOR_5_3_NUM86 (.ZN (XNOR_5_3_NUM86_OUT), .A1 (XNOR_5_1_NUM86_OUT), .A2 (XNOR_5_2_NUM86_OUT));

       wire XNOR_6_1_NUM86_OUT, XNOR_6_2_NUM86_OUT, XNOR_6_3_NUM86_OUT;
       NOR2_X1 XNOR_6_1_NUM86 (.ZN (XNOR_6_1_NUM86_OUT), .A1 (XNOR_3_3_NUM86_OUT), .A2 (GND));
       NOR2_X1 XNOR_6_2_NUM86 (.ZN (XNOR_6_2_NUM86_OUT), .A1 (GND), .A2 (XNOR_4_3_NUM86_OUT));
       NOR2_X1 XNOR_6_3_NUM86 (.ZN (XNOR_6_3_NUM86_OUT), .A1 (XNOR_6_1_NUM86_OUT), .A2 (XNOR_6_2_NUM86_OUT));

       wire XNOR_7_1_NUM86_OUT, XNOR_7_2_NUM86_OUT, XNOR_7_3_NUM86_OUT;
       NOR2_X1 XNOR_7_1_NUM86 (.ZN (XNOR_7_1_NUM86_OUT), .A1 (XNOR_5_3_NUM86_OUT), .A2 (GND));
       NOR2_X1 XNOR_7_2_NUM86 (.ZN (XNOR_7_2_NUM86_OUT), .A1 (GND), .A2 (XNOR_6_3_NUM86_OUT));
       NOR2_X1 XNOR_7_3_NUM86 (.ZN (XNOR_7_3_NUM86_OUT), .A1 (XNOR_7_1_NUM86_OUT), .A2 (XNOR_7_2_NUM86_OUT));

       wire XNOR_8_1_NUM86_OUT, XNOR_8_2_NUM86_OUT, XNOR_8_3_NUM86_OUT;
       NOR2_X1 XNOR_8_1_NUM86 (.ZN (XNOR_8_1_NUM86_OUT), .A1 (XNOR_7_3_NUM86_OUT), .A2 (GND));
       NOR2_X1 XNOR_8_2_NUM86 (.ZN (XNOR_8_2_NUM86_OUT), .A1 (GND), .A2 (N285));
       NOR2_X1 XNOR_8_3_NUM86 (.ZN (N296), .A1 (XNOR_8_1_NUM86_OUT), .A2 (XNOR_8_2_NUM86_OUT));
       NOR2_X1 XNOR_NUM87 (.ZN (N300), .A1 (N263), .A2 (GND));
       NOR2_X1 XNOR_NUM88 (.ZN (N301), .A1 (N288), .A2 (GND));
       NOR2_X1 XNOR_NUM89 (.ZN (N302), .A1 (N289), .A2 (GND));
       NOR2_X1 XNOR_NUM90 (.ZN (N303), .A1 (N290), .A2 (GND));
       NOR2_X1 XNOR_NUM91 (.ZN (N304), .A1 (N291), .A2 (GND));
       NOR2_X1 XNOR_NUM92 (.ZN (N305), .A1 (N292), .A2 (GND));
       NOR2_X1 XNOR_NUM93 (.ZN (N306), .A1 (N293), .A2 (GND));
       NOR2_X1 XNOR_NUM94 (.ZN (N307), .A1 (N294), .A2 (GND));
       NOR2_X1 XNOR_NUM95 (.ZN (N308), .A1 (N295), .A2 (GND));
       NOR2_X1 XNOR_NUM96 (.ZN (N309), .A1 (N296), .A2 (GND));
       NOR2_X1 XNOR_NUM97 (.ZN (N319), .A1 (N296), .A2 (GND));
       NOR2_X1 XNOR_NUM98 (.ZN (N329), .A1 (N296), .A2 (GND));
       wire XNOR_1_1_NUM99_OUT, XNOR_1_2_NUM99_OUT, XNOR_1_3_NUM99_OUT, XNOR_1_4_NUM99_OUT;
       NOR2_X1 XNOR_1_1_NUM99 (.ZN (XNOR_1_1_NUM99_OUT), .A1 (N309), .A2 (GND));
       NOR2_X1 XNOR_1_2_NUM99 (.ZN (XNOR_1_2_NUM99_OUT), .A1 (GND), .A2 (N260));
       NOR2_X1 XNOR_1_3_NUM99 (.ZN (XNOR_1_3_NUM99_OUT), .A1 (XNOR_1_1_NUM99_OUT), .A2 (XNOR_1_2_NUM99_OUT));
       NOR2_X1 XNOR_1_4_NUM99 (.ZN (XNOR_1_4_NUM99_OUT), .A1 (N309), .A2 (N260));
       NOR2_X1 XNOR_1_5_NUM99 (.ZN (N330), .A1 (XNOR_1_3_NUM99_OUT), .A2 (XNOR_1_4_NUM99_OUT));
       wire XNOR_1_1_NUM100_OUT, XNOR_1_2_NUM100_OUT, XNOR_1_3_NUM100_OUT, XNOR_1_4_NUM100_OUT;
       NOR2_X1 XNOR_1_1_NUM100 (.ZN (XNOR_1_1_NUM100_OUT), .A1 (N309), .A2 (GND));
       NOR2_X1 XNOR_1_2_NUM100 (.ZN (XNOR_1_2_NUM100_OUT), .A1 (GND), .A2 (N264));
       NOR2_X1 XNOR_1_3_NUM100 (.ZN (XNOR_1_3_NUM100_OUT), .A1 (XNOR_1_1_NUM100_OUT), .A2 (XNOR_1_2_NUM100_OUT));
       NOR2_X1 XNOR_1_4_NUM100 (.ZN (XNOR_1_4_NUM100_OUT), .A1 (N309), .A2 (N264));
       NOR2_X1 XNOR_1_5_NUM100 (.ZN (N331), .A1 (XNOR_1_3_NUM100_OUT), .A2 (XNOR_1_4_NUM100_OUT));
       wire XNOR_1_1_NUM101_OUT, XNOR_1_2_NUM101_OUT, XNOR_1_3_NUM101_OUT, XNOR_1_4_NUM101_OUT;
       NOR2_X1 XNOR_1_1_NUM101 (.ZN (XNOR_1_1_NUM101_OUT), .A1 (N309), .A2 (GND));
       NOR2_X1 XNOR_1_2_NUM101 (.ZN (XNOR_1_2_NUM101_OUT), .A1 (GND), .A2 (N267));
       NOR2_X1 XNOR_1_3_NUM101 (.ZN (XNOR_1_3_NUM101_OUT), .A1 (XNOR_1_1_NUM101_OUT), .A2 (XNOR_1_2_NUM101_OUT));
       NOR2_X1 XNOR_1_4_NUM101 (.ZN (XNOR_1_4_NUM101_OUT), .A1 (N309), .A2 (N267));
       NOR2_X1 XNOR_1_5_NUM101 (.ZN (N332), .A1 (XNOR_1_3_NUM101_OUT), .A2 (XNOR_1_4_NUM101_OUT));
       wire XNOR_1_1_NUM102_OUT, XNOR_1_2_NUM102_OUT, XNOR_1_3_NUM102_OUT, XNOR_1_4_NUM102_OUT;
       NOR2_X1 XNOR_1_1_NUM102 (.ZN (XNOR_1_1_NUM102_OUT), .A1 (N309), .A2 (GND));
       NOR2_X1 XNOR_1_2_NUM102 (.ZN (XNOR_1_2_NUM102_OUT), .A1 (GND), .A2 (N270));
       NOR2_X1 XNOR_1_3_NUM102 (.ZN (XNOR_1_3_NUM102_OUT), .A1 (XNOR_1_1_NUM102_OUT), .A2 (XNOR_1_2_NUM102_OUT));
       NOR2_X1 XNOR_1_4_NUM102 (.ZN (XNOR_1_4_NUM102_OUT), .A1 (N309), .A2 (N270));
       NOR2_X1 XNOR_1_5_NUM102 (.ZN (N333), .A1 (XNOR_1_3_NUM102_OUT), .A2 (XNOR_1_4_NUM102_OUT));
       wire XNOR_1_1_NUM103_OUT, XNOR_1_2_NUM103_OUT, XNOR_1_3_NUM103_OUT;
       NOR2_X1 XNOR_1_1_NUM103 (.ZN (XNOR_1_1_NUM103_OUT), .A1 (N8), .A2 (GND));
       NOR2_X1 XNOR_1_2_NUM103 (.ZN (XNOR_1_2_NUM103_OUT), .A1 (GND), .A2 (N319));
       NOR2_X1 XNOR_1_3_NUM103 (.ZN (XNOR_1_3_NUM103_OUT), .A1 (XNOR_1_1_NUM103_OUT), .A2 (XNOR_1_2_NUM103_OUT));
       NOR2_X1 XNOR_1_4_NUM103 (.ZN (N334), .A1 (XNOR_1_3_NUM103_OUT), .A2 (GND));
       wire XNOR_1_1_NUM104_OUT, XNOR_1_2_NUM104_OUT, XNOR_1_3_NUM104_OUT, XNOR_1_4_NUM104_OUT;
       NOR2_X1 XNOR_1_1_NUM104 (.ZN (XNOR_1_1_NUM104_OUT), .A1 (N309), .A2 (GND));
       NOR2_X1 XNOR_1_2_NUM104 (.ZN (XNOR_1_2_NUM104_OUT), .A1 (GND), .A2 (N273));
       NOR2_X1 XNOR_1_3_NUM104 (.ZN (XNOR_1_3_NUM104_OUT), .A1 (XNOR_1_1_NUM104_OUT), .A2 (XNOR_1_2_NUM104_OUT));
       NOR2_X1 XNOR_1_4_NUM104 (.ZN (XNOR_1_4_NUM104_OUT), .A1 (N309), .A2 (N273));
       NOR2_X1 XNOR_1_5_NUM104 (.ZN (N335), .A1 (XNOR_1_3_NUM104_OUT), .A2 (XNOR_1_4_NUM104_OUT));
       wire XNOR_1_1_NUM105_OUT, XNOR_1_2_NUM105_OUT, XNOR_1_3_NUM105_OUT;
       NOR2_X1 XNOR_1_1_NUM105 (.ZN (XNOR_1_1_NUM105_OUT), .A1 (N319), .A2 (GND));
       NOR2_X1 XNOR_1_2_NUM105 (.ZN (XNOR_1_2_NUM105_OUT), .A1 (GND), .A2 (N21));
       NOR2_X1 XNOR_1_3_NUM105 (.ZN (XNOR_1_3_NUM105_OUT), .A1 (XNOR_1_1_NUM105_OUT), .A2 (XNOR_1_2_NUM105_OUT));
       NOR2_X1 XNOR_1_4_NUM105 (.ZN (N336), .A1 (XNOR_1_3_NUM105_OUT), .A2 (GND));
       wire XNOR_1_1_NUM106_OUT, XNOR_1_2_NUM106_OUT, XNOR_1_3_NUM106_OUT, XNOR_1_4_NUM106_OUT;
       NOR2_X1 XNOR_1_1_NUM106 (.ZN (XNOR_1_1_NUM106_OUT), .A1 (N309), .A2 (GND));
       NOR2_X1 XNOR_1_2_NUM106 (.ZN (XNOR_1_2_NUM106_OUT), .A1 (GND), .A2 (N276));
       NOR2_X1 XNOR_1_3_NUM106 (.ZN (XNOR_1_3_NUM106_OUT), .A1 (XNOR_1_1_NUM106_OUT), .A2 (XNOR_1_2_NUM106_OUT));
       NOR2_X1 XNOR_1_4_NUM106 (.ZN (XNOR_1_4_NUM106_OUT), .A1 (N309), .A2 (N276));
       NOR2_X1 XNOR_1_5_NUM106 (.ZN (N337), .A1 (XNOR_1_3_NUM106_OUT), .A2 (XNOR_1_4_NUM106_OUT));
       wire XNOR_1_1_NUM107_OUT, XNOR_1_2_NUM107_OUT, XNOR_1_3_NUM107_OUT;
       NOR2_X1 XNOR_1_1_NUM107 (.ZN (XNOR_1_1_NUM107_OUT), .A1 (N319), .A2 (GND));
       NOR2_X1 XNOR_1_2_NUM107 (.ZN (XNOR_1_2_NUM107_OUT), .A1 (GND), .A2 (N34));
       NOR2_X1 XNOR_1_3_NUM107 (.ZN (XNOR_1_3_NUM107_OUT), .A1 (XNOR_1_1_NUM107_OUT), .A2 (XNOR_1_2_NUM107_OUT));
       NOR2_X1 XNOR_1_4_NUM107 (.ZN (N338), .A1 (XNOR_1_3_NUM107_OUT), .A2 (GND));
       wire XNOR_1_1_NUM108_OUT, XNOR_1_2_NUM108_OUT, XNOR_1_3_NUM108_OUT, XNOR_1_4_NUM108_OUT;
       NOR2_X1 XNOR_1_1_NUM108 (.ZN (XNOR_1_1_NUM108_OUT), .A1 (N309), .A2 (GND));
       NOR2_X1 XNOR_1_2_NUM108 (.ZN (XNOR_1_2_NUM108_OUT), .A1 (GND), .A2 (N279));
       NOR2_X1 XNOR_1_3_NUM108 (.ZN (XNOR_1_3_NUM108_OUT), .A1 (XNOR_1_1_NUM108_OUT), .A2 (XNOR_1_2_NUM108_OUT));
       NOR2_X1 XNOR_1_4_NUM108 (.ZN (XNOR_1_4_NUM108_OUT), .A1 (N309), .A2 (N279));
       NOR2_X1 XNOR_1_5_NUM108 (.ZN (N339), .A1 (XNOR_1_3_NUM108_OUT), .A2 (XNOR_1_4_NUM108_OUT));
       wire XNOR_1_1_NUM109_OUT, XNOR_1_2_NUM109_OUT, XNOR_1_3_NUM109_OUT;
       NOR2_X1 XNOR_1_1_NUM109 (.ZN (XNOR_1_1_NUM109_OUT), .A1 (N319), .A2 (GND));
       NOR2_X1 XNOR_1_2_NUM109 (.ZN (XNOR_1_2_NUM109_OUT), .A1 (GND), .A2 (N47));
       NOR2_X1 XNOR_1_3_NUM109 (.ZN (XNOR_1_3_NUM109_OUT), .A1 (XNOR_1_1_NUM109_OUT), .A2 (XNOR_1_2_NUM109_OUT));
       NOR2_X1 XNOR_1_4_NUM109 (.ZN (N340), .A1 (XNOR_1_3_NUM109_OUT), .A2 (GND));
       wire XNOR_1_1_NUM110_OUT, XNOR_1_2_NUM110_OUT, XNOR_1_3_NUM110_OUT, XNOR_1_4_NUM110_OUT;
       NOR2_X1 XNOR_1_1_NUM110 (.ZN (XNOR_1_1_NUM110_OUT), .A1 (N309), .A2 (GND));
       NOR2_X1 XNOR_1_2_NUM110 (.ZN (XNOR_1_2_NUM110_OUT), .A1 (GND), .A2 (N282));
       NOR2_X1 XNOR_1_3_NUM110 (.ZN (XNOR_1_3_NUM110_OUT), .A1 (XNOR_1_1_NUM110_OUT), .A2 (XNOR_1_2_NUM110_OUT));
       NOR2_X1 XNOR_1_4_NUM110 (.ZN (XNOR_1_4_NUM110_OUT), .A1 (N309), .A2 (N282));
       NOR2_X1 XNOR_1_5_NUM110 (.ZN (N341), .A1 (XNOR_1_3_NUM110_OUT), .A2 (XNOR_1_4_NUM110_OUT));
       wire XNOR_1_1_NUM111_OUT, XNOR_1_2_NUM111_OUT, XNOR_1_3_NUM111_OUT;
       NOR2_X1 XNOR_1_1_NUM111 (.ZN (XNOR_1_1_NUM111_OUT), .A1 (N319), .A2 (GND));
       NOR2_X1 XNOR_1_2_NUM111 (.ZN (XNOR_1_2_NUM111_OUT), .A1 (GND), .A2 (N60));
       NOR2_X1 XNOR_1_3_NUM111 (.ZN (XNOR_1_3_NUM111_OUT), .A1 (XNOR_1_1_NUM111_OUT), .A2 (XNOR_1_2_NUM111_OUT));
       NOR2_X1 XNOR_1_4_NUM111 (.ZN (N342), .A1 (XNOR_1_3_NUM111_OUT), .A2 (GND));
       wire XNOR_1_1_NUM112_OUT, XNOR_1_2_NUM112_OUT, XNOR_1_3_NUM112_OUT, XNOR_1_4_NUM112_OUT;
       NOR2_X1 XNOR_1_1_NUM112 (.ZN (XNOR_1_1_NUM112_OUT), .A1 (N309), .A2 (GND));
       NOR2_X1 XNOR_1_2_NUM112 (.ZN (XNOR_1_2_NUM112_OUT), .A1 (GND), .A2 (N285));
       NOR2_X1 XNOR_1_3_NUM112 (.ZN (XNOR_1_3_NUM112_OUT), .A1 (XNOR_1_1_NUM112_OUT), .A2 (XNOR_1_2_NUM112_OUT));
       NOR2_X1 XNOR_1_4_NUM112 (.ZN (XNOR_1_4_NUM112_OUT), .A1 (N309), .A2 (N285));
       NOR2_X1 XNOR_1_5_NUM112 (.ZN (N343), .A1 (XNOR_1_3_NUM112_OUT), .A2 (XNOR_1_4_NUM112_OUT));
       wire XNOR_1_1_NUM113_OUT, XNOR_1_2_NUM113_OUT, XNOR_1_3_NUM113_OUT;
       NOR2_X1 XNOR_1_1_NUM113 (.ZN (XNOR_1_1_NUM113_OUT), .A1 (N319), .A2 (GND));
       NOR2_X1 XNOR_1_2_NUM113 (.ZN (XNOR_1_2_NUM113_OUT), .A1 (GND), .A2 (N73));
       NOR2_X1 XNOR_1_3_NUM113 (.ZN (XNOR_1_3_NUM113_OUT), .A1 (XNOR_1_1_NUM113_OUT), .A2 (XNOR_1_2_NUM113_OUT));
       NOR2_X1 XNOR_1_4_NUM113 (.ZN (N344), .A1 (XNOR_1_3_NUM113_OUT), .A2 (GND));
       wire XNOR_1_1_NUM114_OUT, XNOR_1_2_NUM114_OUT, XNOR_1_3_NUM114_OUT;
       NOR2_X1 XNOR_1_1_NUM114 (.ZN (XNOR_1_1_NUM114_OUT), .A1 (N319), .A2 (GND));
       NOR2_X1 XNOR_1_2_NUM114 (.ZN (XNOR_1_2_NUM114_OUT), .A1 (GND), .A2 (N86));
       NOR2_X1 XNOR_1_3_NUM114 (.ZN (XNOR_1_3_NUM114_OUT), .A1 (XNOR_1_1_NUM114_OUT), .A2 (XNOR_1_2_NUM114_OUT));
       NOR2_X1 XNOR_1_4_NUM114 (.ZN (N345), .A1 (XNOR_1_3_NUM114_OUT), .A2 (GND));
       wire XNOR_1_1_NUM115_OUT, XNOR_1_2_NUM115_OUT, XNOR_1_3_NUM115_OUT;
       NOR2_X1 XNOR_1_1_NUM115 (.ZN (XNOR_1_1_NUM115_OUT), .A1 (N319), .A2 (GND));
       NOR2_X1 XNOR_1_2_NUM115 (.ZN (XNOR_1_2_NUM115_OUT), .A1 (GND), .A2 (N99));
       NOR2_X1 XNOR_1_3_NUM115 (.ZN (XNOR_1_3_NUM115_OUT), .A1 (XNOR_1_1_NUM115_OUT), .A2 (XNOR_1_2_NUM115_OUT));
       NOR2_X1 XNOR_1_4_NUM115 (.ZN (N346), .A1 (XNOR_1_3_NUM115_OUT), .A2 (GND));
       wire XNOR_1_1_NUM116_OUT, XNOR_1_2_NUM116_OUT, XNOR_1_3_NUM116_OUT;
       NOR2_X1 XNOR_1_1_NUM116 (.ZN (XNOR_1_1_NUM116_OUT), .A1 (N319), .A2 (GND));
       NOR2_X1 XNOR_1_2_NUM116 (.ZN (XNOR_1_2_NUM116_OUT), .A1 (GND), .A2 (N112));
       NOR2_X1 XNOR_1_3_NUM116 (.ZN (XNOR_1_3_NUM116_OUT), .A1 (XNOR_1_1_NUM116_OUT), .A2 (XNOR_1_2_NUM116_OUT));
       NOR2_X1 XNOR_1_4_NUM116 (.ZN (N347), .A1 (XNOR_1_3_NUM116_OUT), .A2 (GND));
       wire XNOR_1_1_NUM117_OUT, XNOR_1_2_NUM117_OUT, XNOR_1_3_NUM117_OUT;
       NOR2_X1 XNOR_1_1_NUM117 (.ZN (XNOR_1_1_NUM117_OUT), .A1 (N330), .A2 (GND));
       NOR2_X1 XNOR_1_2_NUM117 (.ZN (XNOR_1_2_NUM117_OUT), .A1 (GND), .A2 (N300));
       NOR2_X1 XNOR_1_3_NUM117 (.ZN (XNOR_1_3_NUM117_OUT), .A1 (XNOR_1_1_NUM117_OUT), .A2 (XNOR_1_2_NUM117_OUT));
       NOR2_X1 XNOR_1_4_NUM117 (.ZN (N348), .A1 (XNOR_1_3_NUM117_OUT), .A2 (GND));
       wire XNOR_1_1_NUM118_OUT, XNOR_1_2_NUM118_OUT, XNOR_1_3_NUM118_OUT;
       NOR2_X1 XNOR_1_1_NUM118 (.ZN (XNOR_1_1_NUM118_OUT), .A1 (N331), .A2 (GND));
       NOR2_X1 XNOR_1_2_NUM118 (.ZN (XNOR_1_2_NUM118_OUT), .A1 (GND), .A2 (N301));
       NOR2_X1 XNOR_1_3_NUM118 (.ZN (XNOR_1_3_NUM118_OUT), .A1 (XNOR_1_1_NUM118_OUT), .A2 (XNOR_1_2_NUM118_OUT));
       NOR2_X1 XNOR_1_4_NUM118 (.ZN (N349), .A1 (XNOR_1_3_NUM118_OUT), .A2 (GND));
       wire XNOR_1_1_NUM119_OUT, XNOR_1_2_NUM119_OUT, XNOR_1_3_NUM119_OUT;
       NOR2_X1 XNOR_1_1_NUM119 (.ZN (XNOR_1_1_NUM119_OUT), .A1 (N332), .A2 (GND));
       NOR2_X1 XNOR_1_2_NUM119 (.ZN (XNOR_1_2_NUM119_OUT), .A1 (GND), .A2 (N302));
       NOR2_X1 XNOR_1_3_NUM119 (.ZN (XNOR_1_3_NUM119_OUT), .A1 (XNOR_1_1_NUM119_OUT), .A2 (XNOR_1_2_NUM119_OUT));
       NOR2_X1 XNOR_1_4_NUM119 (.ZN (N350), .A1 (XNOR_1_3_NUM119_OUT), .A2 (GND));
       wire XNOR_1_1_NUM120_OUT, XNOR_1_2_NUM120_OUT, XNOR_1_3_NUM120_OUT;
       NOR2_X1 XNOR_1_1_NUM120 (.ZN (XNOR_1_1_NUM120_OUT), .A1 (N333), .A2 (GND));
       NOR2_X1 XNOR_1_2_NUM120 (.ZN (XNOR_1_2_NUM120_OUT), .A1 (GND), .A2 (N303));
       NOR2_X1 XNOR_1_3_NUM120 (.ZN (XNOR_1_3_NUM120_OUT), .A1 (XNOR_1_1_NUM120_OUT), .A2 (XNOR_1_2_NUM120_OUT));
       NOR2_X1 XNOR_1_4_NUM120 (.ZN (N351), .A1 (XNOR_1_3_NUM120_OUT), .A2 (GND));
       wire XNOR_1_1_NUM121_OUT, XNOR_1_2_NUM121_OUT, XNOR_1_3_NUM121_OUT;
       NOR2_X1 XNOR_1_1_NUM121 (.ZN (XNOR_1_1_NUM121_OUT), .A1 (N335), .A2 (GND));
       NOR2_X1 XNOR_1_2_NUM121 (.ZN (XNOR_1_2_NUM121_OUT), .A1 (GND), .A2 (N304));
       NOR2_X1 XNOR_1_3_NUM121 (.ZN (XNOR_1_3_NUM121_OUT), .A1 (XNOR_1_1_NUM121_OUT), .A2 (XNOR_1_2_NUM121_OUT));
       NOR2_X1 XNOR_1_4_NUM121 (.ZN (N352), .A1 (XNOR_1_3_NUM121_OUT), .A2 (GND));
       wire XNOR_1_1_NUM122_OUT, XNOR_1_2_NUM122_OUT, XNOR_1_3_NUM122_OUT;
       NOR2_X1 XNOR_1_1_NUM122 (.ZN (XNOR_1_1_NUM122_OUT), .A1 (N337), .A2 (GND));
       NOR2_X1 XNOR_1_2_NUM122 (.ZN (XNOR_1_2_NUM122_OUT), .A1 (GND), .A2 (N305));
       NOR2_X1 XNOR_1_3_NUM122 (.ZN (XNOR_1_3_NUM122_OUT), .A1 (XNOR_1_1_NUM122_OUT), .A2 (XNOR_1_2_NUM122_OUT));
       NOR2_X1 XNOR_1_4_NUM122 (.ZN (N353), .A1 (XNOR_1_3_NUM122_OUT), .A2 (GND));
       wire XNOR_1_1_NUM123_OUT, XNOR_1_2_NUM123_OUT, XNOR_1_3_NUM123_OUT;
       NOR2_X1 XNOR_1_1_NUM123 (.ZN (XNOR_1_1_NUM123_OUT), .A1 (N339), .A2 (GND));
       NOR2_X1 XNOR_1_2_NUM123 (.ZN (XNOR_1_2_NUM123_OUT), .A1 (GND), .A2 (N306));
       NOR2_X1 XNOR_1_3_NUM123 (.ZN (XNOR_1_3_NUM123_OUT), .A1 (XNOR_1_1_NUM123_OUT), .A2 (XNOR_1_2_NUM123_OUT));
       NOR2_X1 XNOR_1_4_NUM123 (.ZN (N354), .A1 (XNOR_1_3_NUM123_OUT), .A2 (GND));
       wire XNOR_1_1_NUM124_OUT, XNOR_1_2_NUM124_OUT, XNOR_1_3_NUM124_OUT;
       NOR2_X1 XNOR_1_1_NUM124 (.ZN (XNOR_1_1_NUM124_OUT), .A1 (N341), .A2 (GND));
       NOR2_X1 XNOR_1_2_NUM124 (.ZN (XNOR_1_2_NUM124_OUT), .A1 (GND), .A2 (N307));
       NOR2_X1 XNOR_1_3_NUM124 (.ZN (XNOR_1_3_NUM124_OUT), .A1 (XNOR_1_1_NUM124_OUT), .A2 (XNOR_1_2_NUM124_OUT));
       NOR2_X1 XNOR_1_4_NUM124 (.ZN (N355), .A1 (XNOR_1_3_NUM124_OUT), .A2 (GND));
       wire XNOR_1_1_NUM125_OUT, XNOR_1_2_NUM125_OUT, XNOR_1_3_NUM125_OUT;
       NOR2_X1 XNOR_1_1_NUM125 (.ZN (XNOR_1_1_NUM125_OUT), .A1 (N343), .A2 (GND));
       NOR2_X1 XNOR_1_2_NUM125 (.ZN (XNOR_1_2_NUM125_OUT), .A1 (GND), .A2 (N308));
       NOR2_X1 XNOR_1_3_NUM125 (.ZN (XNOR_1_3_NUM125_OUT), .A1 (XNOR_1_1_NUM125_OUT), .A2 (XNOR_1_2_NUM125_OUT));
       NOR2_X1 XNOR_1_4_NUM125 (.ZN (N356), .A1 (XNOR_1_3_NUM125_OUT), .A2 (GND));
       wire XNOR_1_1_NUM126_OUT, XNOR_1_2_NUM126_OUT, XNOR_1_3_NUM126_OUT;
       NOR2_X1 XNOR_1_1_NUM126 (.ZN (XNOR_1_1_NUM126_OUT), .A1 (N348), .A2 (GND));
       NOR2_X1 XNOR_1_2_NUM126 (.ZN (XNOR_1_2_NUM126_OUT), .A1 (GND), .A2 (N349));
       NOR2_X1 XNOR_1_3_NUM126 (.ZN (XNOR_1_3_NUM126_OUT), .A1 (XNOR_1_1_NUM126_OUT), .A2 (XNOR_1_2_NUM126_OUT));

       wire XNOR_2_1_NUM126_OUT, XNOR_2_2_NUM126_OUT, XNOR_2_3_NUM126_OUT;
       NOR2_X1 XNOR_2_1_NUM126 (.ZN (XNOR_2_1_NUM126_OUT), .A1 (N350), .A2 (GND));
       NOR2_X1 XNOR_2_2_NUM126 (.ZN (XNOR_2_2_NUM126_OUT), .A1 (GND), .A2 (N351));
       NOR2_X1 XNOR_2_3_NUM126 (.ZN (XNOR_2_3_NUM126_OUT), .A1 (XNOR_2_1_NUM126_OUT), .A2 (XNOR_2_2_NUM126_OUT));

       wire XNOR_3_1_NUM126_OUT, XNOR_3_2_NUM126_OUT, XNOR_3_3_NUM126_OUT;
       NOR2_X1 XNOR_3_1_NUM126 (.ZN (XNOR_3_1_NUM126_OUT), .A1 (N352), .A2 (GND));
       NOR2_X1 XNOR_3_2_NUM126 (.ZN (XNOR_3_2_NUM126_OUT), .A1 (GND), .A2 (N353));
       NOR2_X1 XNOR_3_3_NUM126 (.ZN (XNOR_3_3_NUM126_OUT), .A1 (XNOR_3_1_NUM126_OUT), .A2 (XNOR_3_2_NUM126_OUT));

       wire XNOR_4_1_NUM126_OUT, XNOR_4_2_NUM126_OUT, XNOR_4_3_NUM126_OUT;
       NOR2_X1 XNOR_4_1_NUM126 (.ZN (XNOR_4_1_NUM126_OUT), .A1 (N354), .A2 (GND));
       NOR2_X1 XNOR_4_2_NUM126 (.ZN (XNOR_4_2_NUM126_OUT), .A1 (GND), .A2 (N355));
       NOR2_X1 XNOR_4_3_NUM126 (.ZN (XNOR_4_3_NUM126_OUT), .A1 (XNOR_4_1_NUM126_OUT), .A2 (XNOR_4_2_NUM126_OUT));

       wire XNOR_5_1_NUM126_OUT, XNOR_5_2_NUM126_OUT, XNOR_5_3_NUM126_OUT;
       NOR2_X1 XNOR_5_1_NUM126 (.ZN (XNOR_5_1_NUM126_OUT), .A1 (XNOR_1_3_NUM126_OUT), .A2 (GND));
       NOR2_X1 XNOR_5_2_NUM126 (.ZN (XNOR_5_2_NUM126_OUT), .A1 (GND), .A2 (XNOR_2_3_NUM126_OUT));
       NOR2_X1 XNOR_5_3_NUM126 (.ZN (XNOR_5_3_NUM126_OUT), .A1 (XNOR_5_1_NUM126_OUT), .A2 (XNOR_5_2_NUM126_OUT));

       wire XNOR_6_1_NUM126_OUT, XNOR_6_2_NUM126_OUT, XNOR_6_3_NUM126_OUT;
       NOR2_X1 XNOR_6_1_NUM126 (.ZN (XNOR_6_1_NUM126_OUT), .A1 (XNOR_3_3_NUM126_OUT), .A2 (GND));
       NOR2_X1 XNOR_6_2_NUM126 (.ZN (XNOR_6_2_NUM126_OUT), .A1 (GND), .A2 (XNOR_4_3_NUM126_OUT));
       NOR2_X1 XNOR_6_3_NUM126 (.ZN (XNOR_6_3_NUM126_OUT), .A1 (XNOR_6_1_NUM126_OUT), .A2 (XNOR_6_2_NUM126_OUT));

       wire XNOR_7_1_NUM126_OUT, XNOR_7_2_NUM126_OUT, XNOR_7_3_NUM126_OUT;
       NOR2_X1 XNOR_7_1_NUM126 (.ZN (XNOR_7_1_NUM126_OUT), .A1 (XNOR_5_3_NUM126_OUT), .A2 (GND));
       NOR2_X1 XNOR_7_2_NUM126 (.ZN (XNOR_7_2_NUM126_OUT), .A1 (GND), .A2 (XNOR_6_3_NUM126_OUT));
       NOR2_X1 XNOR_7_3_NUM126 (.ZN (XNOR_7_3_NUM126_OUT), .A1 (XNOR_7_1_NUM126_OUT), .A2 (XNOR_7_2_NUM126_OUT));

       wire XNOR_8_1_NUM126_OUT, XNOR_8_2_NUM126_OUT, XNOR_8_3_NUM126_OUT;
       NOR2_X1 XNOR_8_1_NUM126 (.ZN (XNOR_8_1_NUM126_OUT), .A1 (XNOR_7_3_NUM126_OUT), .A2 (GND));
       NOR2_X1 XNOR_8_2_NUM126 (.ZN (XNOR_8_2_NUM126_OUT), .A1 (GND), .A2 (N356));
       NOR2_X1 XNOR_8_3_NUM126 (.ZN (N357), .A1 (XNOR_8_1_NUM126_OUT), .A2 (XNOR_8_2_NUM126_OUT));
       NOR2_X1 XNOR_NUM127 (.ZN (N360), .A1 (N357), .A2 (GND));
       NOR2_X1 XNOR_NUM128 (.ZN (N370), .A1 (N357), .A2 (GND));
       wire XNOR_1_1_NUM129_OUT, XNOR_1_2_NUM129_OUT, XNOR_1_3_NUM129_OUT;
       NOR2_X1 XNOR_1_1_NUM129 (.ZN (XNOR_1_1_NUM129_OUT), .A1 (N14), .A2 (GND));
       NOR2_X1 XNOR_1_2_NUM129 (.ZN (XNOR_1_2_NUM129_OUT), .A1 (GND), .A2 (N360));
       NOR2_X1 XNOR_1_3_NUM129 (.ZN (XNOR_1_3_NUM129_OUT), .A1 (XNOR_1_1_NUM129_OUT), .A2 (XNOR_1_2_NUM129_OUT));
       NOR2_X1 XNOR_1_4_NUM129 (.ZN (N371), .A1 (XNOR_1_3_NUM129_OUT), .A2 (GND));
       wire XNOR_1_1_NUM130_OUT, XNOR_1_2_NUM130_OUT, XNOR_1_3_NUM130_OUT;
       NOR2_X1 XNOR_1_1_NUM130 (.ZN (XNOR_1_1_NUM130_OUT), .A1 (N360), .A2 (GND));
       NOR2_X1 XNOR_1_2_NUM130 (.ZN (XNOR_1_2_NUM130_OUT), .A1 (GND), .A2 (N27));
       NOR2_X1 XNOR_1_3_NUM130 (.ZN (XNOR_1_3_NUM130_OUT), .A1 (XNOR_1_1_NUM130_OUT), .A2 (XNOR_1_2_NUM130_OUT));
       NOR2_X1 XNOR_1_4_NUM130 (.ZN (N372), .A1 (XNOR_1_3_NUM130_OUT), .A2 (GND));
       wire XNOR_1_1_NUM131_OUT, XNOR_1_2_NUM131_OUT, XNOR_1_3_NUM131_OUT;
       NOR2_X1 XNOR_1_1_NUM131 (.ZN (XNOR_1_1_NUM131_OUT), .A1 (N360), .A2 (GND));
       NOR2_X1 XNOR_1_2_NUM131 (.ZN (XNOR_1_2_NUM131_OUT), .A1 (GND), .A2 (N40));
       NOR2_X1 XNOR_1_3_NUM131 (.ZN (XNOR_1_3_NUM131_OUT), .A1 (XNOR_1_1_NUM131_OUT), .A2 (XNOR_1_2_NUM131_OUT));
       NOR2_X1 XNOR_1_4_NUM131 (.ZN (N373), .A1 (XNOR_1_3_NUM131_OUT), .A2 (GND));
       wire XNOR_1_1_NUM132_OUT, XNOR_1_2_NUM132_OUT, XNOR_1_3_NUM132_OUT;
       NOR2_X1 XNOR_1_1_NUM132 (.ZN (XNOR_1_1_NUM132_OUT), .A1 (N360), .A2 (GND));
       NOR2_X1 XNOR_1_2_NUM132 (.ZN (XNOR_1_2_NUM132_OUT), .A1 (GND), .A2 (N53));
       NOR2_X1 XNOR_1_3_NUM132 (.ZN (XNOR_1_3_NUM132_OUT), .A1 (XNOR_1_1_NUM132_OUT), .A2 (XNOR_1_2_NUM132_OUT));
       NOR2_X1 XNOR_1_4_NUM132 (.ZN (N374), .A1 (XNOR_1_3_NUM132_OUT), .A2 (GND));
       wire XNOR_1_1_NUM133_OUT, XNOR_1_2_NUM133_OUT, XNOR_1_3_NUM133_OUT;
       NOR2_X1 XNOR_1_1_NUM133 (.ZN (XNOR_1_1_NUM133_OUT), .A1 (N360), .A2 (GND));
       NOR2_X1 XNOR_1_2_NUM133 (.ZN (XNOR_1_2_NUM133_OUT), .A1 (GND), .A2 (N66));
       NOR2_X1 XNOR_1_3_NUM133 (.ZN (XNOR_1_3_NUM133_OUT), .A1 (XNOR_1_1_NUM133_OUT), .A2 (XNOR_1_2_NUM133_OUT));
       NOR2_X1 XNOR_1_4_NUM133 (.ZN (N375), .A1 (XNOR_1_3_NUM133_OUT), .A2 (GND));
       wire XNOR_1_1_NUM134_OUT, XNOR_1_2_NUM134_OUT, XNOR_1_3_NUM134_OUT;
       NOR2_X1 XNOR_1_1_NUM134 (.ZN (XNOR_1_1_NUM134_OUT), .A1 (N360), .A2 (GND));
       NOR2_X1 XNOR_1_2_NUM134 (.ZN (XNOR_1_2_NUM134_OUT), .A1 (GND), .A2 (N79));
       NOR2_X1 XNOR_1_3_NUM134 (.ZN (XNOR_1_3_NUM134_OUT), .A1 (XNOR_1_1_NUM134_OUT), .A2 (XNOR_1_2_NUM134_OUT));
       NOR2_X1 XNOR_1_4_NUM134 (.ZN (N376), .A1 (XNOR_1_3_NUM134_OUT), .A2 (GND));
       wire XNOR_1_1_NUM135_OUT, XNOR_1_2_NUM135_OUT, XNOR_1_3_NUM135_OUT;
       NOR2_X1 XNOR_1_1_NUM135 (.ZN (XNOR_1_1_NUM135_OUT), .A1 (N360), .A2 (GND));
       NOR2_X1 XNOR_1_2_NUM135 (.ZN (XNOR_1_2_NUM135_OUT), .A1 (GND), .A2 (N92));
       NOR2_X1 XNOR_1_3_NUM135 (.ZN (XNOR_1_3_NUM135_OUT), .A1 (XNOR_1_1_NUM135_OUT), .A2 (XNOR_1_2_NUM135_OUT));
       NOR2_X1 XNOR_1_4_NUM135 (.ZN (N377), .A1 (XNOR_1_3_NUM135_OUT), .A2 (GND));
       wire XNOR_1_1_NUM136_OUT, XNOR_1_2_NUM136_OUT, XNOR_1_3_NUM136_OUT;
       NOR2_X1 XNOR_1_1_NUM136 (.ZN (XNOR_1_1_NUM136_OUT), .A1 (N360), .A2 (GND));
       NOR2_X1 XNOR_1_2_NUM136 (.ZN (XNOR_1_2_NUM136_OUT), .A1 (GND), .A2 (N105));
       NOR2_X1 XNOR_1_3_NUM136 (.ZN (XNOR_1_3_NUM136_OUT), .A1 (XNOR_1_1_NUM136_OUT), .A2 (XNOR_1_2_NUM136_OUT));
       NOR2_X1 XNOR_1_4_NUM136 (.ZN (N378), .A1 (XNOR_1_3_NUM136_OUT), .A2 (GND));
       wire XNOR_1_1_NUM137_OUT, XNOR_1_2_NUM137_OUT, XNOR_1_3_NUM137_OUT;
       NOR2_X1 XNOR_1_1_NUM137 (.ZN (XNOR_1_1_NUM137_OUT), .A1 (N360), .A2 (GND));
       NOR2_X1 XNOR_1_2_NUM137 (.ZN (XNOR_1_2_NUM137_OUT), .A1 (GND), .A2 (N115));
       NOR2_X1 XNOR_1_3_NUM137 (.ZN (XNOR_1_3_NUM137_OUT), .A1 (XNOR_1_1_NUM137_OUT), .A2 (XNOR_1_2_NUM137_OUT));
       NOR2_X1 XNOR_1_4_NUM137 (.ZN (N379), .A1 (XNOR_1_3_NUM137_OUT), .A2 (GND));
       wire XNOR_1_1_NUM138_OUT, XNOR_1_2_NUM138_OUT, XNOR_1_3_NUM138_OUT;
       NOR2_X1 XNOR_1_1_NUM138 (.ZN (XNOR_1_1_NUM138_OUT), .A1 (N4), .A2 (GND));
       NOR2_X1 XNOR_1_2_NUM138 (.ZN (XNOR_1_2_NUM138_OUT), .A1 (GND), .A2 (N242));
       NOR2_X1 XNOR_1_3_NUM138 (.ZN (XNOR_1_3_NUM138_OUT), .A1 (XNOR_1_1_NUM138_OUT), .A2 (XNOR_1_2_NUM138_OUT));

       wire XNOR_2_1_NUM138_OUT, XNOR_2_2_NUM138_OUT, XNOR_2_3_NUM138_OUT;
       NOR2_X1 XNOR_2_1_NUM138 (.ZN (XNOR_2_1_NUM138_OUT), .A1 (N334), .A2 (GND));
       NOR2_X1 XNOR_2_2_NUM138 (.ZN (XNOR_2_2_NUM138_OUT), .A1 (GND), .A2 (N371));
       NOR2_X1 XNOR_2_3_NUM138 (.ZN (XNOR_2_3_NUM138_OUT), .A1 (XNOR_2_1_NUM138_OUT), .A2 (XNOR_2_2_NUM138_OUT));

       wire XNOR_3_1_NUM138_OUT, XNOR_3_2_NUM138_OUT, XNOR_3_3_NUM138_OUT;
       NOR2_X1 XNOR_3_1_NUM138 (.ZN (XNOR_3_1_NUM138_OUT), .A1 (XNOR_1_3_NUM138_OUT), .A2 (GND));
       NOR2_X1 XNOR_3_2_NUM138 (.ZN (XNOR_3_2_NUM138_OUT), .A1 (GND), .A2 (XNOR_2_3_NUM138_OUT));
       NOR2_X1 XNOR_3_3_NUM138 (.ZN (XNOR_3_3_NUM138_OUT), .A1 (XNOR_3_1_NUM138_OUT), .A2 (XNOR_3_2_NUM138_OUT));

       NOR2_X1 XNOR_4_1_NUM138 (.ZN (N380), .A1 (XNOR_3_3_NUM138_OUT), .A2 (GND));
       wire XNOR_1_1_NUM139_OUT, XNOR_1_2_NUM139_OUT, XNOR_1_3_NUM139_OUT;
       NOR2_X1 XNOR_1_1_NUM139 (.ZN (XNOR_1_1_NUM139_OUT), .A1 (N246), .A2 (GND));
       NOR2_X1 XNOR_1_2_NUM139 (.ZN (XNOR_1_2_NUM139_OUT), .A1 (GND), .A2 (N336));
       NOR2_X1 XNOR_1_3_NUM139 (.ZN (XNOR_1_3_NUM139_OUT), .A1 (XNOR_1_1_NUM139_OUT), .A2 (XNOR_1_2_NUM139_OUT));

       wire XNOR_2_1_NUM139_OUT, XNOR_2_2_NUM139_OUT, XNOR_2_3_NUM139_OUT;
       NOR2_X1 XNOR_2_1_NUM139 (.ZN (XNOR_2_1_NUM139_OUT), .A1 (N372), .A2 (GND));
       NOR2_X1 XNOR_2_2_NUM139 (.ZN (XNOR_2_2_NUM139_OUT), .A1 (GND), .A2 (N17));
       NOR2_X1 XNOR_2_3_NUM139 (.ZN (XNOR_2_3_NUM139_OUT), .A1 (XNOR_2_1_NUM139_OUT), .A2 (XNOR_2_2_NUM139_OUT));

       wire XNOR_3_1_NUM139_OUT, XNOR_3_2_NUM139_OUT, XNOR_3_3_NUM139_OUT;
       NOR2_X1 XNOR_3_1_NUM139 (.ZN (XNOR_3_1_NUM139_OUT), .A1 (XNOR_1_3_NUM139_OUT), .A2 (GND));
       NOR2_X1 XNOR_3_2_NUM139 (.ZN (XNOR_3_2_NUM139_OUT), .A1 (GND), .A2 (XNOR_2_3_NUM139_OUT));
       NOR2_X1 XNOR_3_3_NUM139 (.ZN (XNOR_3_3_NUM139_OUT), .A1 (XNOR_3_1_NUM139_OUT), .A2 (XNOR_3_2_NUM139_OUT));

       NOR2_X1 XNOR_4_1_NUM139 (.ZN (N381), .A1 (XNOR_3_3_NUM139_OUT), .A2 (GND));
       wire XNOR_1_1_NUM140_OUT, XNOR_1_2_NUM140_OUT, XNOR_1_3_NUM140_OUT;
       NOR2_X1 XNOR_1_1_NUM140 (.ZN (XNOR_1_1_NUM140_OUT), .A1 (N250), .A2 (GND));
       NOR2_X1 XNOR_1_2_NUM140 (.ZN (XNOR_1_2_NUM140_OUT), .A1 (GND), .A2 (N338));
       NOR2_X1 XNOR_1_3_NUM140 (.ZN (XNOR_1_3_NUM140_OUT), .A1 (XNOR_1_1_NUM140_OUT), .A2 (XNOR_1_2_NUM140_OUT));

       wire XNOR_2_1_NUM140_OUT, XNOR_2_2_NUM140_OUT, XNOR_2_3_NUM140_OUT;
       NOR2_X1 XNOR_2_1_NUM140 (.ZN (XNOR_2_1_NUM140_OUT), .A1 (N373), .A2 (GND));
       NOR2_X1 XNOR_2_2_NUM140 (.ZN (XNOR_2_2_NUM140_OUT), .A1 (GND), .A2 (N30));
       NOR2_X1 XNOR_2_3_NUM140 (.ZN (XNOR_2_3_NUM140_OUT), .A1 (XNOR_2_1_NUM140_OUT), .A2 (XNOR_2_2_NUM140_OUT));

       wire XNOR_3_1_NUM140_OUT, XNOR_3_2_NUM140_OUT, XNOR_3_3_NUM140_OUT;
       NOR2_X1 XNOR_3_1_NUM140 (.ZN (XNOR_3_1_NUM140_OUT), .A1 (XNOR_1_3_NUM140_OUT), .A2 (GND));
       NOR2_X1 XNOR_3_2_NUM140 (.ZN (XNOR_3_2_NUM140_OUT), .A1 (GND), .A2 (XNOR_2_3_NUM140_OUT));
       NOR2_X1 XNOR_3_3_NUM140 (.ZN (XNOR_3_3_NUM140_OUT), .A1 (XNOR_3_1_NUM140_OUT), .A2 (XNOR_3_2_NUM140_OUT));

       NOR2_X1 XNOR_4_1_NUM140 (.ZN (N386), .A1 (XNOR_3_3_NUM140_OUT), .A2 (GND));
       wire XNOR_1_1_NUM141_OUT, XNOR_1_2_NUM141_OUT, XNOR_1_3_NUM141_OUT;
       NOR2_X1 XNOR_1_1_NUM141 (.ZN (XNOR_1_1_NUM141_OUT), .A1 (N254), .A2 (GND));
       NOR2_X1 XNOR_1_2_NUM141 (.ZN (XNOR_1_2_NUM141_OUT), .A1 (GND), .A2 (N340));
       NOR2_X1 XNOR_1_3_NUM141 (.ZN (XNOR_1_3_NUM141_OUT), .A1 (XNOR_1_1_NUM141_OUT), .A2 (XNOR_1_2_NUM141_OUT));

       wire XNOR_2_1_NUM141_OUT, XNOR_2_2_NUM141_OUT, XNOR_2_3_NUM141_OUT;
       NOR2_X1 XNOR_2_1_NUM141 (.ZN (XNOR_2_1_NUM141_OUT), .A1 (N374), .A2 (GND));
       NOR2_X1 XNOR_2_2_NUM141 (.ZN (XNOR_2_2_NUM141_OUT), .A1 (GND), .A2 (N43));
       NOR2_X1 XNOR_2_3_NUM141 (.ZN (XNOR_2_3_NUM141_OUT), .A1 (XNOR_2_1_NUM141_OUT), .A2 (XNOR_2_2_NUM141_OUT));

       wire XNOR_3_1_NUM141_OUT, XNOR_3_2_NUM141_OUT, XNOR_3_3_NUM141_OUT;
       NOR2_X1 XNOR_3_1_NUM141 (.ZN (XNOR_3_1_NUM141_OUT), .A1 (XNOR_1_3_NUM141_OUT), .A2 (GND));
       NOR2_X1 XNOR_3_2_NUM141 (.ZN (XNOR_3_2_NUM141_OUT), .A1 (GND), .A2 (XNOR_2_3_NUM141_OUT));
       NOR2_X1 XNOR_3_3_NUM141 (.ZN (XNOR_3_3_NUM141_OUT), .A1 (XNOR_3_1_NUM141_OUT), .A2 (XNOR_3_2_NUM141_OUT));

       NOR2_X1 XNOR_4_1_NUM141 (.ZN (N393), .A1 (XNOR_3_3_NUM141_OUT), .A2 (GND));
       wire XNOR_1_1_NUM142_OUT, XNOR_1_2_NUM142_OUT, XNOR_1_3_NUM142_OUT;
       NOR2_X1 XNOR_1_1_NUM142 (.ZN (XNOR_1_1_NUM142_OUT), .A1 (N255), .A2 (GND));
       NOR2_X1 XNOR_1_2_NUM142 (.ZN (XNOR_1_2_NUM142_OUT), .A1 (GND), .A2 (N342));
       NOR2_X1 XNOR_1_3_NUM142 (.ZN (XNOR_1_3_NUM142_OUT), .A1 (XNOR_1_1_NUM142_OUT), .A2 (XNOR_1_2_NUM142_OUT));

       wire XNOR_2_1_NUM142_OUT, XNOR_2_2_NUM142_OUT, XNOR_2_3_NUM142_OUT;
       NOR2_X1 XNOR_2_1_NUM142 (.ZN (XNOR_2_1_NUM142_OUT), .A1 (N375), .A2 (GND));
       NOR2_X1 XNOR_2_2_NUM142 (.ZN (XNOR_2_2_NUM142_OUT), .A1 (GND), .A2 (N56));
       NOR2_X1 XNOR_2_3_NUM142 (.ZN (XNOR_2_3_NUM142_OUT), .A1 (XNOR_2_1_NUM142_OUT), .A2 (XNOR_2_2_NUM142_OUT));

       wire XNOR_3_1_NUM142_OUT, XNOR_3_2_NUM142_OUT, XNOR_3_3_NUM142_OUT;
       NOR2_X1 XNOR_3_1_NUM142 (.ZN (XNOR_3_1_NUM142_OUT), .A1 (XNOR_1_3_NUM142_OUT), .A2 (GND));
       NOR2_X1 XNOR_3_2_NUM142 (.ZN (XNOR_3_2_NUM142_OUT), .A1 (GND), .A2 (XNOR_2_3_NUM142_OUT));
       NOR2_X1 XNOR_3_3_NUM142 (.ZN (XNOR_3_3_NUM142_OUT), .A1 (XNOR_3_1_NUM142_OUT), .A2 (XNOR_3_2_NUM142_OUT));

       NOR2_X1 XNOR_4_1_NUM142 (.ZN (N399), .A1 (XNOR_3_3_NUM142_OUT), .A2 (GND));
       wire XNOR_1_1_NUM143_OUT, XNOR_1_2_NUM143_OUT, XNOR_1_3_NUM143_OUT;
       NOR2_X1 XNOR_1_1_NUM143 (.ZN (XNOR_1_1_NUM143_OUT), .A1 (N256), .A2 (GND));
       NOR2_X1 XNOR_1_2_NUM143 (.ZN (XNOR_1_2_NUM143_OUT), .A1 (GND), .A2 (N344));
       NOR2_X1 XNOR_1_3_NUM143 (.ZN (XNOR_1_3_NUM143_OUT), .A1 (XNOR_1_1_NUM143_OUT), .A2 (XNOR_1_2_NUM143_OUT));

       wire XNOR_2_1_NUM143_OUT, XNOR_2_2_NUM143_OUT, XNOR_2_3_NUM143_OUT;
       NOR2_X1 XNOR_2_1_NUM143 (.ZN (XNOR_2_1_NUM143_OUT), .A1 (N376), .A2 (GND));
       NOR2_X1 XNOR_2_2_NUM143 (.ZN (XNOR_2_2_NUM143_OUT), .A1 (GND), .A2 (N69));
       NOR2_X1 XNOR_2_3_NUM143 (.ZN (XNOR_2_3_NUM143_OUT), .A1 (XNOR_2_1_NUM143_OUT), .A2 (XNOR_2_2_NUM143_OUT));

       wire XNOR_3_1_NUM143_OUT, XNOR_3_2_NUM143_OUT, XNOR_3_3_NUM143_OUT;
       NOR2_X1 XNOR_3_1_NUM143 (.ZN (XNOR_3_1_NUM143_OUT), .A1 (XNOR_1_3_NUM143_OUT), .A2 (GND));
       NOR2_X1 XNOR_3_2_NUM143 (.ZN (XNOR_3_2_NUM143_OUT), .A1 (GND), .A2 (XNOR_2_3_NUM143_OUT));
       NOR2_X1 XNOR_3_3_NUM143 (.ZN (XNOR_3_3_NUM143_OUT), .A1 (XNOR_3_1_NUM143_OUT), .A2 (XNOR_3_2_NUM143_OUT));

       NOR2_X1 XNOR_4_1_NUM143 (.ZN (N404), .A1 (XNOR_3_3_NUM143_OUT), .A2 (GND));
       wire XNOR_1_1_NUM144_OUT, XNOR_1_2_NUM144_OUT, XNOR_1_3_NUM144_OUT;
       NOR2_X1 XNOR_1_1_NUM144 (.ZN (XNOR_1_1_NUM144_OUT), .A1 (N257), .A2 (GND));
       NOR2_X1 XNOR_1_2_NUM144 (.ZN (XNOR_1_2_NUM144_OUT), .A1 (GND), .A2 (N345));
       NOR2_X1 XNOR_1_3_NUM144 (.ZN (XNOR_1_3_NUM144_OUT), .A1 (XNOR_1_1_NUM144_OUT), .A2 (XNOR_1_2_NUM144_OUT));

       wire XNOR_2_1_NUM144_OUT, XNOR_2_2_NUM144_OUT, XNOR_2_3_NUM144_OUT;
       NOR2_X1 XNOR_2_1_NUM144 (.ZN (XNOR_2_1_NUM144_OUT), .A1 (N377), .A2 (GND));
       NOR2_X1 XNOR_2_2_NUM144 (.ZN (XNOR_2_2_NUM144_OUT), .A1 (GND), .A2 (N82));
       NOR2_X1 XNOR_2_3_NUM144 (.ZN (XNOR_2_3_NUM144_OUT), .A1 (XNOR_2_1_NUM144_OUT), .A2 (XNOR_2_2_NUM144_OUT));

       wire XNOR_3_1_NUM144_OUT, XNOR_3_2_NUM144_OUT, XNOR_3_3_NUM144_OUT;
       NOR2_X1 XNOR_3_1_NUM144 (.ZN (XNOR_3_1_NUM144_OUT), .A1 (XNOR_1_3_NUM144_OUT), .A2 (GND));
       NOR2_X1 XNOR_3_2_NUM144 (.ZN (XNOR_3_2_NUM144_OUT), .A1 (GND), .A2 (XNOR_2_3_NUM144_OUT));
       NOR2_X1 XNOR_3_3_NUM144 (.ZN (XNOR_3_3_NUM144_OUT), .A1 (XNOR_3_1_NUM144_OUT), .A2 (XNOR_3_2_NUM144_OUT));

       NOR2_X1 XNOR_4_1_NUM144 (.ZN (N407), .A1 (XNOR_3_3_NUM144_OUT), .A2 (GND));
       wire XNOR_1_1_NUM145_OUT, XNOR_1_2_NUM145_OUT, XNOR_1_3_NUM145_OUT;
       NOR2_X1 XNOR_1_1_NUM145 (.ZN (XNOR_1_1_NUM145_OUT), .A1 (N258), .A2 (GND));
       NOR2_X1 XNOR_1_2_NUM145 (.ZN (XNOR_1_2_NUM145_OUT), .A1 (GND), .A2 (N346));
       NOR2_X1 XNOR_1_3_NUM145 (.ZN (XNOR_1_3_NUM145_OUT), .A1 (XNOR_1_1_NUM145_OUT), .A2 (XNOR_1_2_NUM145_OUT));

       wire XNOR_2_1_NUM145_OUT, XNOR_2_2_NUM145_OUT, XNOR_2_3_NUM145_OUT;
       NOR2_X1 XNOR_2_1_NUM145 (.ZN (XNOR_2_1_NUM145_OUT), .A1 (N378), .A2 (GND));
       NOR2_X1 XNOR_2_2_NUM145 (.ZN (XNOR_2_2_NUM145_OUT), .A1 (GND), .A2 (N95));
       NOR2_X1 XNOR_2_3_NUM145 (.ZN (XNOR_2_3_NUM145_OUT), .A1 (XNOR_2_1_NUM145_OUT), .A2 (XNOR_2_2_NUM145_OUT));

       wire XNOR_3_1_NUM145_OUT, XNOR_3_2_NUM145_OUT, XNOR_3_3_NUM145_OUT;
       NOR2_X1 XNOR_3_1_NUM145 (.ZN (XNOR_3_1_NUM145_OUT), .A1 (XNOR_1_3_NUM145_OUT), .A2 (GND));
       NOR2_X1 XNOR_3_2_NUM145 (.ZN (XNOR_3_2_NUM145_OUT), .A1 (GND), .A2 (XNOR_2_3_NUM145_OUT));
       NOR2_X1 XNOR_3_3_NUM145 (.ZN (XNOR_3_3_NUM145_OUT), .A1 (XNOR_3_1_NUM145_OUT), .A2 (XNOR_3_2_NUM145_OUT));

       NOR2_X1 XNOR_4_1_NUM145 (.ZN (N411), .A1 (XNOR_3_3_NUM145_OUT), .A2 (GND));
       wire XNOR_1_1_NUM146_OUT, XNOR_1_2_NUM146_OUT, XNOR_1_3_NUM146_OUT;
       NOR2_X1 XNOR_1_1_NUM146 (.ZN (XNOR_1_1_NUM146_OUT), .A1 (N259), .A2 (GND));
       NOR2_X1 XNOR_1_2_NUM146 (.ZN (XNOR_1_2_NUM146_OUT), .A1 (GND), .A2 (N347));
       NOR2_X1 XNOR_1_3_NUM146 (.ZN (XNOR_1_3_NUM146_OUT), .A1 (XNOR_1_1_NUM146_OUT), .A2 (XNOR_1_2_NUM146_OUT));

       wire XNOR_2_1_NUM146_OUT, XNOR_2_2_NUM146_OUT, XNOR_2_3_NUM146_OUT;
       NOR2_X1 XNOR_2_1_NUM146 (.ZN (XNOR_2_1_NUM146_OUT), .A1 (N379), .A2 (GND));
       NOR2_X1 XNOR_2_2_NUM146 (.ZN (XNOR_2_2_NUM146_OUT), .A1 (GND), .A2 (N108));
       NOR2_X1 XNOR_2_3_NUM146 (.ZN (XNOR_2_3_NUM146_OUT), .A1 (XNOR_2_1_NUM146_OUT), .A2 (XNOR_2_2_NUM146_OUT));

       wire XNOR_3_1_NUM146_OUT, XNOR_3_2_NUM146_OUT, XNOR_3_3_NUM146_OUT;
       NOR2_X1 XNOR_3_1_NUM146 (.ZN (XNOR_3_1_NUM146_OUT), .A1 (XNOR_1_3_NUM146_OUT), .A2 (GND));
       NOR2_X1 XNOR_3_2_NUM146 (.ZN (XNOR_3_2_NUM146_OUT), .A1 (GND), .A2 (XNOR_2_3_NUM146_OUT));
       NOR2_X1 XNOR_3_3_NUM146 (.ZN (XNOR_3_3_NUM146_OUT), .A1 (XNOR_3_1_NUM146_OUT), .A2 (XNOR_3_2_NUM146_OUT));

       NOR2_X1 XNOR_4_1_NUM146 (.ZN (N414), .A1 (XNOR_3_3_NUM146_OUT), .A2 (GND));
       NOR2_X1 XNOR_NUM147 (.ZN (N415), .A1 (N380), .A2 (GND));
       wire XNOR_1_1_NUM148_OUT, XNOR_1_2_NUM148_OUT, XNOR_1_3_NUM148_OUT;
       NOR2_X1 XNOR_1_1_NUM148 (.ZN (XNOR_1_1_NUM148_OUT), .A1 (N381), .A2 (GND));
       NOR2_X1 XNOR_1_2_NUM148 (.ZN (XNOR_1_2_NUM148_OUT), .A1 (GND), .A2 (N386));
       NOR2_X1 XNOR_1_3_NUM148 (.ZN (XNOR_1_3_NUM148_OUT), .A1 (XNOR_1_1_NUM148_OUT), .A2 (XNOR_1_2_NUM148_OUT));

       wire XNOR_2_1_NUM148_OUT, XNOR_2_2_NUM148_OUT, XNOR_2_3_NUM148_OUT;
       NOR2_X1 XNOR_2_1_NUM148 (.ZN (XNOR_2_1_NUM148_OUT), .A1 (N393), .A2 (GND));
       NOR2_X1 XNOR_2_2_NUM148 (.ZN (XNOR_2_2_NUM148_OUT), .A1 (GND), .A2 (N399));
       NOR2_X1 XNOR_2_3_NUM148 (.ZN (XNOR_2_3_NUM148_OUT), .A1 (XNOR_2_1_NUM148_OUT), .A2 (XNOR_2_2_NUM148_OUT));

       wire XNOR_3_1_NUM148_OUT, XNOR_3_2_NUM148_OUT, XNOR_3_3_NUM148_OUT;
       NOR2_X1 XNOR_3_1_NUM148 (.ZN (XNOR_3_1_NUM148_OUT), .A1 (N404), .A2 (GND));
       NOR2_X1 XNOR_3_2_NUM148 (.ZN (XNOR_3_2_NUM148_OUT), .A1 (GND), .A2 (N407));
       NOR2_X1 XNOR_3_3_NUM148 (.ZN (XNOR_3_3_NUM148_OUT), .A1 (XNOR_3_1_NUM148_OUT), .A2 (XNOR_3_2_NUM148_OUT));

       wire XNOR_4_1_NUM148_OUT, XNOR_4_2_NUM148_OUT, XNOR_4_3_NUM148_OUT;
       NOR2_X1 XNOR_4_1_NUM148 (.ZN (XNOR_4_1_NUM148_OUT), .A1 (N411), .A2 (GND));
       NOR2_X1 XNOR_4_2_NUM148 (.ZN (XNOR_4_2_NUM148_OUT), .A1 (GND), .A2 (N414));
       NOR2_X1 XNOR_4_3_NUM148 (.ZN (XNOR_4_3_NUM148_OUT), .A1 (XNOR_4_1_NUM148_OUT), .A2 (XNOR_4_2_NUM148_OUT));

       wire XNOR_5_1_NUM148_OUT, XNOR_5_2_NUM148_OUT, XNOR_5_3_NUM148_OUT;
       NOR2_X1 XNOR_5_1_NUM148 (.ZN (XNOR_5_1_NUM148_OUT), .A1 (XNOR_1_3_NUM148_OUT), .A2 (GND));
       NOR2_X1 XNOR_5_2_NUM148 (.ZN (XNOR_5_2_NUM148_OUT), .A1 (GND), .A2 (XNOR_2_3_NUM148_OUT));
       NOR2_X1 XNOR_5_3_NUM148 (.ZN (XNOR_5_3_NUM148_OUT), .A1 (XNOR_5_1_NUM148_OUT), .A2 (XNOR_5_2_NUM148_OUT));

       wire XNOR_6_1_NUM148_OUT, XNOR_6_2_NUM148_OUT, XNOR_6_3_NUM148_OUT;
       NOR2_X1 XNOR_6_1_NUM148 (.ZN (XNOR_6_1_NUM148_OUT), .A1 (XNOR_3_3_NUM148_OUT), .A2 (GND));
       NOR2_X1 XNOR_6_2_NUM148 (.ZN (XNOR_6_2_NUM148_OUT), .A1 (GND), .A2 (XNOR_4_3_NUM148_OUT));
       NOR2_X1 XNOR_6_3_NUM148 (.ZN (XNOR_6_3_NUM148_OUT), .A1 (XNOR_6_1_NUM148_OUT), .A2 (XNOR_6_2_NUM148_OUT));

       wire XNOR_7_1_NUM148_OUT, XNOR_7_2_NUM148_OUT;
       NOR2_X1 XNOR_7_1_NUM148 (.ZN (XNOR_7_1_NUM148_OUT), .A1 (XNOR_5_3_NUM148_OUT), .A2 (GND));
       NOR2_X1 XNOR_7_2_NUM148 (.ZN (XNOR_7_2_NUM148_OUT), .A1 (GND), .A2 (XNOR_6_3_NUM148_OUT));
       NOR2_X1 XNOR_7_3_NUM148 (.ZN (N416), .A1 (XNOR_7_1_NUM148_OUT), .A2 (XNOR_7_2_NUM148_OUT));
       NOR2_X1 XNOR_NUM149 (.ZN (N417), .A1 (N393), .A2 (GND));
       NOR2_X1 XNOR_NUM150 (.ZN (N418), .A1 (N404), .A2 (GND));
       NOR2_X1 XNOR_NUM151 (.ZN (N419), .A1 (N407), .A2 (GND));
       NOR2_X1 XNOR_NUM152 (.ZN (N420), .A1 (N411), .A2 (GND));
       NOR2_X1 XNOR_NUM153 (.ZN (N421), .A1 (N415), .A2 (N416));
       wire XNOR_1_1_NUM154_OUT, XNOR_1_2_NUM154_OUT, XNOR_1_3_NUM154_OUT;
       NOR2_X1 XNOR_1_1_NUM154 (.ZN (XNOR_1_1_NUM154_OUT), .A1 (N386), .A2 (GND));
       NOR2_X1 XNOR_1_2_NUM154 (.ZN (XNOR_1_2_NUM154_OUT), .A1 (GND), .A2 (N417));
       NOR2_X1 XNOR_1_3_NUM154 (.ZN (XNOR_1_3_NUM154_OUT), .A1 (XNOR_1_1_NUM154_OUT), .A2 (XNOR_1_2_NUM154_OUT));
       NOR2_X1 XNOR_1_4_NUM154 (.ZN (N422), .A1 (XNOR_1_3_NUM154_OUT), .A2 (GND));
       wire XNOR_1_1_NUM155_OUT, XNOR_1_2_NUM155_OUT, XNOR_1_3_NUM155_OUT;
       NOR2_X1 XNOR_1_1_NUM155 (.ZN (XNOR_1_1_NUM155_OUT), .A1 (N386), .A2 (GND));
       NOR2_X1 XNOR_1_2_NUM155 (.ZN (XNOR_1_2_NUM155_OUT), .A1 (GND), .A2 (N393));
       NOR2_X1 XNOR_1_3_NUM155 (.ZN (XNOR_1_3_NUM155_OUT), .A1 (XNOR_1_1_NUM155_OUT), .A2 (XNOR_1_2_NUM155_OUT));

       wire XNOR_2_1_NUM155_OUT, XNOR_2_2_NUM155_OUT, XNOR_2_3_NUM155_OUT;
       NOR2_X1 XNOR_2_1_NUM155 (.ZN (XNOR_2_1_NUM155_OUT), .A1 (N418), .A2 (GND));
       NOR2_X1 XNOR_2_2_NUM155 (.ZN (XNOR_2_2_NUM155_OUT), .A1 (GND), .A2 (N399));
       NOR2_X1 XNOR_2_3_NUM155 (.ZN (XNOR_2_3_NUM155_OUT), .A1 (XNOR_2_1_NUM155_OUT), .A2 (XNOR_2_2_NUM155_OUT));

       wire XNOR_3_1_NUM155_OUT, XNOR_3_2_NUM155_OUT, XNOR_3_3_NUM155_OUT;
       NOR2_X1 XNOR_3_1_NUM155 (.ZN (XNOR_3_1_NUM155_OUT), .A1 (XNOR_1_3_NUM155_OUT), .A2 (GND));
       NOR2_X1 XNOR_3_2_NUM155 (.ZN (XNOR_3_2_NUM155_OUT), .A1 (GND), .A2 (XNOR_2_3_NUM155_OUT));
       NOR2_X1 XNOR_3_3_NUM155 (.ZN (XNOR_3_3_NUM155_OUT), .A1 (XNOR_3_1_NUM155_OUT), .A2 (XNOR_3_2_NUM155_OUT));

       NOR2_X1 XNOR_4_1_NUM155 (.ZN (N425), .A1 (XNOR_3_3_NUM155_OUT), .A2 (GND));
       wire XNOR_1_1_NUM156_OUT, XNOR_1_2_NUM156_OUT, XNOR_1_3_NUM156_OUT;
       NOR2_X1 XNOR_1_1_NUM156 (.ZN (XNOR_1_1_NUM156_OUT), .A1 (N399), .A2 (GND));
       NOR2_X1 XNOR_1_2_NUM156 (.ZN (XNOR_1_2_NUM156_OUT), .A1 (GND), .A2 (N393));
       NOR2_X1 XNOR_1_3_NUM156 (.ZN (XNOR_1_3_NUM156_OUT), .A1 (XNOR_1_1_NUM156_OUT), .A2 (XNOR_1_2_NUM156_OUT));

       wire XNOR_2_1_NUM156_OUT, XNOR_2_2_NUM156_OUT, XNOR_2_3_NUM156_OUT;
       NOR2_X1 XNOR_2_1_NUM156 (.ZN (XNOR_2_1_NUM156_OUT), .A1 (N419), .A2 (GND));
       NOR2_X1 XNOR_2_2_NUM156 (.ZN (XNOR_2_2_NUM156_OUT), .A1 (GND), .A2 (XNOR_1_3_NUM156_OUT));
       NOR2_X1 XNOR_2_3_NUM156 (.ZN (XNOR_2_3_NUM156_OUT), .A1 (XNOR_2_1_NUM156_OUT), .A2 (XNOR_2_2_NUM156_OUT));

       NOR2_X1 XNOR_3_1_NUM156 (.ZN (N428), .A1 (XNOR_2_3_NUM156_OUT), .A2 (GND));
       wire XNOR_1_1_NUM157_OUT, XNOR_1_2_NUM157_OUT, XNOR_1_3_NUM157_OUT;
       NOR2_X1 XNOR_1_1_NUM157 (.ZN (XNOR_1_1_NUM157_OUT), .A1 (N386), .A2 (GND));
       NOR2_X1 XNOR_1_2_NUM157 (.ZN (XNOR_1_2_NUM157_OUT), .A1 (GND), .A2 (N393));
       NOR2_X1 XNOR_1_3_NUM157 (.ZN (XNOR_1_3_NUM157_OUT), .A1 (XNOR_1_1_NUM157_OUT), .A2 (XNOR_1_2_NUM157_OUT));

       wire XNOR_2_1_NUM157_OUT, XNOR_2_2_NUM157_OUT, XNOR_2_3_NUM157_OUT;
       NOR2_X1 XNOR_2_1_NUM157 (.ZN (XNOR_2_1_NUM157_OUT), .A1 (N407), .A2 (GND));
       NOR2_X1 XNOR_2_2_NUM157 (.ZN (XNOR_2_2_NUM157_OUT), .A1 (GND), .A2 (N420));
       NOR2_X1 XNOR_2_3_NUM157 (.ZN (XNOR_2_3_NUM157_OUT), .A1 (XNOR_2_1_NUM157_OUT), .A2 (XNOR_2_2_NUM157_OUT));

       wire XNOR_3_1_NUM157_OUT, XNOR_3_2_NUM157_OUT, XNOR_3_3_NUM157_OUT;
       NOR2_X1 XNOR_3_1_NUM157 (.ZN (XNOR_3_1_NUM157_OUT), .A1 (XNOR_1_3_NUM157_OUT), .A2 (GND));
       NOR2_X1 XNOR_3_2_NUM157 (.ZN (XNOR_3_2_NUM157_OUT), .A1 (GND), .A2 (XNOR_2_3_NUM157_OUT));
       NOR2_X1 XNOR_3_3_NUM157 (.ZN (XNOR_3_3_NUM157_OUT), .A1 (XNOR_3_1_NUM157_OUT), .A2 (XNOR_3_2_NUM157_OUT));

       NOR2_X1 XNOR_4_1_NUM157 (.ZN (N429), .A1 (XNOR_3_3_NUM157_OUT), .A2 (GND));
       wire XNOR_1_1_NUM158_OUT, XNOR_1_2_NUM158_OUT, XNOR_1_3_NUM158_OUT;
       NOR2_X1 XNOR_1_1_NUM158 (.ZN (XNOR_1_1_NUM158_OUT), .A1 (N381), .A2 (GND));
       NOR2_X1 XNOR_1_2_NUM158 (.ZN (XNOR_1_2_NUM158_OUT), .A1 (GND), .A2 (N386));
       NOR2_X1 XNOR_1_3_NUM158 (.ZN (XNOR_1_3_NUM158_OUT), .A1 (XNOR_1_1_NUM158_OUT), .A2 (XNOR_1_2_NUM158_OUT));

       wire XNOR_2_1_NUM158_OUT, XNOR_2_2_NUM158_OUT, XNOR_2_3_NUM158_OUT;
       NOR2_X1 XNOR_2_1_NUM158 (.ZN (XNOR_2_1_NUM158_OUT), .A1 (N422), .A2 (GND));
       NOR2_X1 XNOR_2_2_NUM158 (.ZN (XNOR_2_2_NUM158_OUT), .A1 (GND), .A2 (N399));
       NOR2_X1 XNOR_2_3_NUM158 (.ZN (XNOR_2_3_NUM158_OUT), .A1 (XNOR_2_1_NUM158_OUT), .A2 (XNOR_2_2_NUM158_OUT));

       wire XNOR_3_1_NUM158_OUT, XNOR_3_2_NUM158_OUT, XNOR_3_3_NUM158_OUT;
       NOR2_X1 XNOR_3_1_NUM158 (.ZN (XNOR_3_1_NUM158_OUT), .A1 (XNOR_1_3_NUM158_OUT), .A2 (GND));
       NOR2_X1 XNOR_3_2_NUM158 (.ZN (XNOR_3_2_NUM158_OUT), .A1 (GND), .A2 (XNOR_2_3_NUM158_OUT));
       NOR2_X1 XNOR_3_3_NUM158 (.ZN (XNOR_3_3_NUM158_OUT), .A1 (XNOR_3_1_NUM158_OUT), .A2 (XNOR_3_2_NUM158_OUT));

       NOR2_X1 XNOR_4_1_NUM158 (.ZN (N430), .A1 (XNOR_3_3_NUM158_OUT), .A2 (GND));
       wire XNOR_1_1_NUM159_OUT, XNOR_1_2_NUM159_OUT, XNOR_1_3_NUM159_OUT;
       NOR2_X1 XNOR_1_1_NUM159 (.ZN (XNOR_1_1_NUM159_OUT), .A1 (N381), .A2 (GND));
       NOR2_X1 XNOR_1_2_NUM159 (.ZN (XNOR_1_2_NUM159_OUT), .A1 (GND), .A2 (N386));
       NOR2_X1 XNOR_1_3_NUM159 (.ZN (XNOR_1_3_NUM159_OUT), .A1 (XNOR_1_1_NUM159_OUT), .A2 (XNOR_1_2_NUM159_OUT));

       wire XNOR_2_1_NUM159_OUT, XNOR_2_2_NUM159_OUT, XNOR_2_3_NUM159_OUT;
       NOR2_X1 XNOR_2_1_NUM159 (.ZN (XNOR_2_1_NUM159_OUT), .A1 (N425), .A2 (GND));
       NOR2_X1 XNOR_2_2_NUM159 (.ZN (XNOR_2_2_NUM159_OUT), .A1 (GND), .A2 (N428));
       NOR2_X1 XNOR_2_3_NUM159 (.ZN (XNOR_2_3_NUM159_OUT), .A1 (XNOR_2_1_NUM159_OUT), .A2 (XNOR_2_2_NUM159_OUT));

       wire XNOR_3_1_NUM159_OUT, XNOR_3_2_NUM159_OUT, XNOR_3_3_NUM159_OUT;
       NOR2_X1 XNOR_3_1_NUM159 (.ZN (XNOR_3_1_NUM159_OUT), .A1 (XNOR_1_3_NUM159_OUT), .A2 (GND));
       NOR2_X1 XNOR_3_2_NUM159 (.ZN (XNOR_3_2_NUM159_OUT), .A1 (GND), .A2 (XNOR_2_3_NUM159_OUT));
       NOR2_X1 XNOR_3_3_NUM159 (.ZN (XNOR_3_3_NUM159_OUT), .A1 (XNOR_3_1_NUM159_OUT), .A2 (XNOR_3_2_NUM159_OUT));

       NOR2_X1 XNOR_4_1_NUM159 (.ZN (N431), .A1 (XNOR_3_3_NUM159_OUT), .A2 (GND));
       wire XNOR_1_1_NUM160_OUT, XNOR_1_2_NUM160_OUT, XNOR_1_3_NUM160_OUT;
       NOR2_X1 XNOR_1_1_NUM160 (.ZN (XNOR_1_1_NUM160_OUT), .A1 (N381), .A2 (GND));
       NOR2_X1 XNOR_1_2_NUM160 (.ZN (XNOR_1_2_NUM160_OUT), .A1 (GND), .A2 (N422));
       NOR2_X1 XNOR_1_3_NUM160 (.ZN (XNOR_1_3_NUM160_OUT), .A1 (XNOR_1_1_NUM160_OUT), .A2 (XNOR_1_2_NUM160_OUT));

       wire XNOR_2_1_NUM160_OUT, XNOR_2_2_NUM160_OUT, XNOR_2_3_NUM160_OUT;
       NOR2_X1 XNOR_2_1_NUM160 (.ZN (XNOR_2_1_NUM160_OUT), .A1 (N425), .A2 (GND));
       NOR2_X1 XNOR_2_2_NUM160 (.ZN (XNOR_2_2_NUM160_OUT), .A1 (GND), .A2 (N429));
       NOR2_X1 XNOR_2_3_NUM160 (.ZN (XNOR_2_3_NUM160_OUT), .A1 (XNOR_2_1_NUM160_OUT), .A2 (XNOR_2_2_NUM160_OUT));

       wire XNOR_3_1_NUM160_OUT, XNOR_3_2_NUM160_OUT, XNOR_3_3_NUM160_OUT;
       NOR2_X1 XNOR_3_1_NUM160 (.ZN (XNOR_3_1_NUM160_OUT), .A1 (XNOR_1_3_NUM160_OUT), .A2 (GND));
       NOR2_X1 XNOR_3_2_NUM160 (.ZN (XNOR_3_2_NUM160_OUT), .A1 (GND), .A2 (XNOR_2_3_NUM160_OUT));
       NOR2_X1 XNOR_3_3_NUM160 (.ZN (XNOR_3_3_NUM160_OUT), .A1 (XNOR_3_1_NUM160_OUT), .A2 (XNOR_3_2_NUM160_OUT));

       NOR2_X1 XNOR_4_1_NUM160 (.ZN (N432), .A1 (XNOR_3_3_NUM160_OUT), .A2 (GND));


       wire XNOR_1_1_N223_TERMINATION_OUT, XNOR_1_2_N223_TERMINATION_OUT;
       NOR2_X1 XNOR_1_1_N223_TERMINATION (.ZN (XNOR_1_1_N223_TERMINATION_OUT), .A1 (N223), .A2 (GND));
       NOR2_X1 XNOR_1_2_N223_TERMINATION (.ZN (N223_TERMINATION), .A1 (XNOR_1_1_N223_TERMINATION_OUT), .A2 (XNOR_1_2_N223_TERMINATION_OUT));

       wire XNOR_1_1_N329_TERMINATION_OUT, XNOR_1_2_N329_TERMINATION_OUT;
       NOR2_X1 XNOR_1_1_N329_TERMINATION (.ZN (XNOR_1_1_N329_TERMINATION_OUT), .A1 (N329), .A2 (GND));
       NOR2_X1 XNOR_1_2_N329_TERMINATION (.ZN (N329_TERMINATION), .A1 (XNOR_1_1_N329_TERMINATION_OUT), .A2 (XNOR_1_2_N329_TERMINATION_OUT));

       wire XNOR_1_1_N370_TERMINATION_OUT, XNOR_1_2_N370_TERMINATION_OUT;
       NOR2_X1 XNOR_1_1_N370_TERMINATION (.ZN (XNOR_1_1_N370_TERMINATION_OUT), .A1 (N370), .A2 (GND));
       NOR2_X1 XNOR_1_2_N370_TERMINATION (.ZN (N370_TERMINATION), .A1 (XNOR_1_1_N370_TERMINATION_OUT), .A2 (XNOR_1_2_N370_TERMINATION_OUT));

       wire XNOR_1_1_N421_TERMINATION_OUT, XNOR_1_2_N421_TERMINATION_OUT;
       NOR2_X1 XNOR_1_1_N421_TERMINATION (.ZN (XNOR_1_1_N421_TERMINATION_OUT), .A1 (N421), .A2 (GND));
       NOR2_X1 XNOR_1_2_N421_TERMINATION (.ZN (N421_TERMINATION), .A1 (XNOR_1_1_N421_TERMINATION_OUT), .A2 (XNOR_1_2_N421_TERMINATION_OUT));

       wire XNOR_1_1_N430_TERMINATION_OUT, XNOR_1_2_N430_TERMINATION_OUT;
       NOR2_X1 XNOR_1_1_N430_TERMINATION (.ZN (XNOR_1_1_N430_TERMINATION_OUT), .A1 (N430), .A2 (GND));
       NOR2_X1 XNOR_1_2_N430_TERMINATION (.ZN (N430_TERMINATION), .A1 (XNOR_1_1_N430_TERMINATION_OUT), .A2 (XNOR_1_2_N430_TERMINATION_OUT));

       wire XNOR_1_1_N431_TERMINATION_OUT, XNOR_1_2_N431_TERMINATION_OUT;
       NOR2_X1 XNOR_1_1_N431_TERMINATION (.ZN (XNOR_1_1_N431_TERMINATION_OUT), .A1 (N431), .A2 (GND));
       NOR2_X1 XNOR_1_2_N431_TERMINATION (.ZN (N431_TERMINATION), .A1 (XNOR_1_1_N431_TERMINATION_OUT), .A2 (XNOR_1_2_N431_TERMINATION_OUT));

       wire XNOR_1_1_N432_TERMINATION_OUT, XNOR_1_2_N432_TERMINATION_OUT;
       NOR2_X1 XNOR_1_1_N432_TERMINATION (.ZN (XNOR_1_1_N432_TERMINATION_OUT), .A1 (N432), .A2 (GND));
       NOR2_X1 XNOR_1_2_N432_TERMINATION (.ZN (N432_TERMINATION), .A1 (XNOR_1_1_N432_TERMINATION_OUT), .A2 (XNOR_1_2_N432_TERMINATION_OUT));


endmodule
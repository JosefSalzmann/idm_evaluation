* circuit: nor inv chain with alternating nor inputs
simulator lang=spice

*.PARAM pw=<sed>pw<sed>as
.PARAM supp=0.8V slope=0.1fs
.PARAM t_init0=0.1ns t_init1=0.174ns
.PARAM baseVal=0V peakVal=0.8V tend=1.0ns


.LIB /home/s11777724/involution_tool_library_files/backend/spice/fet.inc CMG

* main circuit
.INCLUDE /home/s11777724/involution_tool_library_files/backend/spice/cell/NOR2_X1.sp

**** SPECTRE Back Annotation
.option spef='/home/s11777724/JS/idm_evaluation/nor_inv_chain_altered_inputs_b/place_and_route/nor_inv_chain_altered_inputs_b_generic_parasitics.spef'
****

.TEMP 25
.OPTION
+ INGOLD=2
+ PARHIER=LOCAL
*+ POST=CSDF
+ PROBE
+ BRIEF
+ ACCURATE
+ ABSVAR=0.0001
+ DVDT=2
+ RELTOL=1e-11
*+ DELMAX=100fs
+ dc_pivot_check=yes

* vdd
VDD VDD GND 0.8v

VIN myin GND PWL 0ns baseVal t_init0 baseVal 't_init0+slope' peakVal t_init1 peakVal 't_init1+slope' baseVal

* circuit under test
XNOR0 GND myin STAGE0 VDD VDD GND GND NOR2_X1
XNOR2 GND STAGE0 STAGE2 VDD VDD GND GND NOR2_X1
XNOR3 GND STAGE2 STAGE3 VDD VDD GND GND NOR2_X1
XNOR4 GND STAGE3 STAGE4 VDD VDD GND GND NOR2_X1
XNOR5 GND STAGE4 STAGE5 VDD VDD GND GND NOR2_X1
XNOR6 GND STAGE5 STAGE6 VDD VDD GND GND NOR2_X1
XNOR7 GND STAGE6 STAGE7 VDD VDD GND GND NOR2_X1
XNOR8 GND STAGE7 STAGE8 VDD VDD GND GND NOR2_X1
XNOR9 GND STAGE8 STAGE9 VDD VDD GND GND NOR2_X1
XNOR10 GND STAGE9 STAGE10 VDD VDD GND GND NOR2_X1
XNOR11 STAGE10 GND STAGE11 VDD VDD GND GND NOR2_X1
XNOR12 GND STAGE11 STAGE12 VDD VDD GND GND NOR2_X1
XNOR13 STAGE12 GND STAGE13 VDD VDD GND GND NOR2_X1
XNOR14 GND STAGE13 STAGE14 VDD VDD GND GND NOR2_X1
XNOR15 STAGE14 GND STAGE15 VDD VDD GND GND NOR2_X1
XNOR16 GND STAGE15 STAGE16 VDD VDD GND GND NOR2_X1
XNOR17 STAGE16 GND STAGE17 VDD VDD GND GND NOR2_X1
XNOR18 GND STAGE17 STAGE18 VDD VDD GND GND NOR2_X1
XNOR19 STAGE18 GND STAGE19 VDD VDD GND GND NOR2_X1
XNOR20 GND STAGE19 STAGE20 VDD VDD GND GND NOR2_X1
XNOR21 STAGE20 GND STAGE21 VDD VDD GND GND NOR2_X1
XNOR22 GND STAGE21 STAGE22 VDD VDD GND GND NOR2_X1
XNOR23 STAGE22 GND STAGE23 VDD VDD GND GND NOR2_X1
XNOR24 GND STAGE23 STAGE24 VDD VDD GND GND NOR2_X1
XNOR25 STAGE24 GND myout VDD VDD GND GND NOR2_X1
C_TERM myout GND 0.0779pF

.PROBE TRAN V(STAGE9) V(STAGE10)
+ V(STAGE11) V(STAGE12) V(STAGE13) V(STAGE14) V(STAGE15)
+ V(STAGE16) V(STAGE17) V(STAGE18) V(STAGE19) V(STAGE20)
+ V(STAGE21)
.TRAN 0.1ps tend
.END

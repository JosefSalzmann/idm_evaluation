module c6288_NOR_template (N1_PWL,N18_PWL,N35_PWL,N52_PWL,N69_PWL,N86_PWL,N103_PWL,N120_PWL,N137_PWL,N154_PWL,N171_PWL,
            N188_PWL,N205_PWL,N222_PWL,N239_PWL,N256_PWL,N273_PWL,N290_PWL,N307_PWL,N324_PWL,N341_PWL,N358_PWL,
            N375_PWL,N392_PWL,N409_PWL,N426_PWL,N443_PWL,N460_PWL,N477_PWL,N494_PWL,N511_PWL,N528_PWL,
            N545_TERMINATION,N1581_TERMINATION,N1901_TERMINATION,N2223_TERMINATION,N2548_TERMINATION,
            N2877_TERMINATION,N3211_TERMINATION,N3552_TERMINATION,N3895_TERMINATION,N4241_TERMINATION,
            N4591_TERMINATION,N4946_TERMINATION,N5308_TERMINATION,N5672_TERMINATION,N5971_TERMINATION,
            N6123_TERMINATION,N6150_TERMINATION,N6160_TERMINATION,N6170_TERMINATION,N6180_TERMINATION,
            N6190_TERMINATION,N6200_TERMINATION,N6210_TERMINATION,N6220_TERMINATION,N6230_TERMINATION,
            N6240_TERMINATION,N6250_TERMINATION,N6260_TERMINATION,N6270_TERMINATION,N6280_TERMINATION,
            N6287_TERMINATION,N6288_TERMINATION);

      input N1_PWL,N18_PWL,N35_PWL,N52_PWL,N69_PWL,N86_PWL,N103_PWL,N120_PWL,N137_PWL,N154_PWL,N171_PWL,
            N188_PWL,N205_PWL,N222_PWL,N239_PWL,N256_PWL,N273_PWL,N290_PWL,N307_PWL,N324_PWL,N341_PWL,N358_PWL,
            N375_PWL,N392_PWL,N409_PWL,N426_PWL,N443_PWL,N460_PWL,N477_PWL,N494_PWL,N511_PWL,N528_PWL;

      output N545_TERMINATION,N1581_TERMINATION,N1901_TERMINATION,N2223_TERMINATION,N2548_TERMINATION,
            N2877_TERMINATION,N3211_TERMINATION,N3552_TERMINATION,N3895_TERMINATION,N4241_TERMINATION,
            N4591_TERMINATION,N4946_TERMINATION,N5308_TERMINATION,N5672_TERMINATION,N5971_TERMINATION,
            N6123_TERMINATION,N6150_TERMINATION,N6160_TERMINATION,N6170_TERMINATION,N6180_TERMINATION,
            N6190_TERMINATION,N6200_TERMINATION,N6210_TERMINATION,N6220_TERMINATION,N6230_TERMINATION,
            N6240_TERMINATION,N6250_TERMINATION,N6260_TERMINATION,N6270_TERMINATION,N6280_TERMINATION,
            N6287_TERMINATION,N6288_TERMINATION;

      wire GND = 1'b0;
      wire XNOR_1_1_N1_PULSESHAPING_OUT, XNOR_1_2_N1_PULSESHAPING_OUT, XNOR_1_3_N1_PULSESHAPING_OUT, XNOR_1_4_N1_PULSESHAPING_OUT, XNOR_1_5_N1_PULSESHAPING_OUT, XNOR_1_6_N1_PULSESHAPING_OUT;
      NOR2_X1 XNOR_1_1_N1_PULSESHAPING (.ZN (XNOR_1_1_N1_PULSESHAPING_OUT), .A1 (N1_PWL), .A2 (GND));
      NOR2_X1 XNOR_1_2_N1_PULSESHAPING (.ZN (XNOR_1_2_N1_PULSESHAPING_OUT), .A1 (XNOR_1_1_N1_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_3_N1_PULSESHAPING (.ZN (XNOR_1_3_N1_PULSESHAPING_OUT), .A1 (XNOR_1_2_N1_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_4_N1_PULSESHAPING (.ZN (XNOR_1_4_N1_PULSESHAPING_OUT), .A1 (XNOR_1_3_N1_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_5_N1_PULSESHAPING (.ZN (XNOR_1_5_N1_PULSESHAPING_OUT), .A1 (XNOR_1_4_N1_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_6_N1_PULSESHAPING (.ZN (XNOR_1_6_N1_PULSESHAPING_OUT), .A1 (XNOR_1_5_N1_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_7_N1_PULSESHAPING (.ZN (N1), .A1 (XNOR_1_6_N1_PULSESHAPING_OUT), .A2 (GND));

      wire XNOR_1_1_N18_PULSESHAPING_OUT, XNOR_1_2_N18_PULSESHAPING_OUT, XNOR_1_3_N18_PULSESHAPING_OUT, XNOR_1_4_N18_PULSESHAPING_OUT, XNOR_1_5_N18_PULSESHAPING_OUT, XNOR_1_6_N18_PULSESHAPING_OUT;
      NOR2_X1 XNOR_1_1_N18_PULSESHAPING (.ZN (XNOR_1_1_N18_PULSESHAPING_OUT), .A1 (N18_PWL), .A2 (GND));
      NOR2_X1 XNOR_1_2_N18_PULSESHAPING (.ZN (XNOR_1_2_N18_PULSESHAPING_OUT), .A1 (XNOR_1_1_N18_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_3_N18_PULSESHAPING (.ZN (XNOR_1_3_N18_PULSESHAPING_OUT), .A1 (XNOR_1_2_N18_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_4_N18_PULSESHAPING (.ZN (XNOR_1_4_N18_PULSESHAPING_OUT), .A1 (XNOR_1_3_N18_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_5_N18_PULSESHAPING (.ZN (XNOR_1_5_N18_PULSESHAPING_OUT), .A1 (XNOR_1_4_N18_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_6_N18_PULSESHAPING (.ZN (XNOR_1_6_N18_PULSESHAPING_OUT), .A1 (XNOR_1_5_N18_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_7_N18_PULSESHAPING (.ZN (N18), .A1 (XNOR_1_6_N18_PULSESHAPING_OUT), .A2 (GND));

      wire XNOR_1_1_N35_PULSESHAPING_OUT, XNOR_1_2_N35_PULSESHAPING_OUT, XNOR_1_3_N35_PULSESHAPING_OUT, XNOR_1_4_N35_PULSESHAPING_OUT, XNOR_1_5_N35_PULSESHAPING_OUT, XNOR_1_6_N35_PULSESHAPING_OUT;
      NOR2_X1 XNOR_1_1_N35_PULSESHAPING (.ZN (XNOR_1_1_N35_PULSESHAPING_OUT), .A1 (N35_PWL), .A2 (GND));
      NOR2_X1 XNOR_1_2_N35_PULSESHAPING (.ZN (XNOR_1_2_N35_PULSESHAPING_OUT), .A1 (XNOR_1_1_N35_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_3_N35_PULSESHAPING (.ZN (XNOR_1_3_N35_PULSESHAPING_OUT), .A1 (XNOR_1_2_N35_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_4_N35_PULSESHAPING (.ZN (XNOR_1_4_N35_PULSESHAPING_OUT), .A1 (XNOR_1_3_N35_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_5_N35_PULSESHAPING (.ZN (XNOR_1_5_N35_PULSESHAPING_OUT), .A1 (XNOR_1_4_N35_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_6_N35_PULSESHAPING (.ZN (XNOR_1_6_N35_PULSESHAPING_OUT), .A1 (XNOR_1_5_N35_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_7_N35_PULSESHAPING (.ZN (N35), .A1 (XNOR_1_6_N35_PULSESHAPING_OUT), .A2 (GND));

      wire XNOR_1_1_N52_PULSESHAPING_OUT, XNOR_1_2_N52_PULSESHAPING_OUT, XNOR_1_3_N52_PULSESHAPING_OUT, XNOR_1_4_N52_PULSESHAPING_OUT, XNOR_1_5_N52_PULSESHAPING_OUT, XNOR_1_6_N52_PULSESHAPING_OUT;
      NOR2_X1 XNOR_1_1_N52_PULSESHAPING (.ZN (XNOR_1_1_N52_PULSESHAPING_OUT), .A1 (N52_PWL), .A2 (GND));
      NOR2_X1 XNOR_1_2_N52_PULSESHAPING (.ZN (XNOR_1_2_N52_PULSESHAPING_OUT), .A1 (XNOR_1_1_N52_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_3_N52_PULSESHAPING (.ZN (XNOR_1_3_N52_PULSESHAPING_OUT), .A1 (XNOR_1_2_N52_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_4_N52_PULSESHAPING (.ZN (XNOR_1_4_N52_PULSESHAPING_OUT), .A1 (XNOR_1_3_N52_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_5_N52_PULSESHAPING (.ZN (XNOR_1_5_N52_PULSESHAPING_OUT), .A1 (XNOR_1_4_N52_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_6_N52_PULSESHAPING (.ZN (XNOR_1_6_N52_PULSESHAPING_OUT), .A1 (XNOR_1_5_N52_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_7_N52_PULSESHAPING (.ZN (N52), .A1 (XNOR_1_6_N52_PULSESHAPING_OUT), .A2 (GND));

      wire XNOR_1_1_N69_PULSESHAPING_OUT, XNOR_1_2_N69_PULSESHAPING_OUT, XNOR_1_3_N69_PULSESHAPING_OUT, XNOR_1_4_N69_PULSESHAPING_OUT, XNOR_1_5_N69_PULSESHAPING_OUT, XNOR_1_6_N69_PULSESHAPING_OUT;
      NOR2_X1 XNOR_1_1_N69_PULSESHAPING (.ZN (XNOR_1_1_N69_PULSESHAPING_OUT), .A1 (N69_PWL), .A2 (GND));
      NOR2_X1 XNOR_1_2_N69_PULSESHAPING (.ZN (XNOR_1_2_N69_PULSESHAPING_OUT), .A1 (XNOR_1_1_N69_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_3_N69_PULSESHAPING (.ZN (XNOR_1_3_N69_PULSESHAPING_OUT), .A1 (XNOR_1_2_N69_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_4_N69_PULSESHAPING (.ZN (XNOR_1_4_N69_PULSESHAPING_OUT), .A1 (XNOR_1_3_N69_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_5_N69_PULSESHAPING (.ZN (XNOR_1_5_N69_PULSESHAPING_OUT), .A1 (XNOR_1_4_N69_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_6_N69_PULSESHAPING (.ZN (XNOR_1_6_N69_PULSESHAPING_OUT), .A1 (XNOR_1_5_N69_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_7_N69_PULSESHAPING (.ZN (N69), .A1 (XNOR_1_6_N69_PULSESHAPING_OUT), .A2 (GND));

      wire XNOR_1_1_N86_PULSESHAPING_OUT, XNOR_1_2_N86_PULSESHAPING_OUT, XNOR_1_3_N86_PULSESHAPING_OUT, XNOR_1_4_N86_PULSESHAPING_OUT, XNOR_1_5_N86_PULSESHAPING_OUT, XNOR_1_6_N86_PULSESHAPING_OUT;
      NOR2_X1 XNOR_1_1_N86_PULSESHAPING (.ZN (XNOR_1_1_N86_PULSESHAPING_OUT), .A1 (N86_PWL), .A2 (GND));
      NOR2_X1 XNOR_1_2_N86_PULSESHAPING (.ZN (XNOR_1_2_N86_PULSESHAPING_OUT), .A1 (XNOR_1_1_N86_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_3_N86_PULSESHAPING (.ZN (XNOR_1_3_N86_PULSESHAPING_OUT), .A1 (XNOR_1_2_N86_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_4_N86_PULSESHAPING (.ZN (XNOR_1_4_N86_PULSESHAPING_OUT), .A1 (XNOR_1_3_N86_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_5_N86_PULSESHAPING (.ZN (XNOR_1_5_N86_PULSESHAPING_OUT), .A1 (XNOR_1_4_N86_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_6_N86_PULSESHAPING (.ZN (XNOR_1_6_N86_PULSESHAPING_OUT), .A1 (XNOR_1_5_N86_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_7_N86_PULSESHAPING (.ZN (N86), .A1 (XNOR_1_6_N86_PULSESHAPING_OUT), .A2 (GND));

      wire XNOR_1_1_N103_PULSESHAPING_OUT, XNOR_1_2_N103_PULSESHAPING_OUT, XNOR_1_3_N103_PULSESHAPING_OUT, XNOR_1_4_N103_PULSESHAPING_OUT, XNOR_1_5_N103_PULSESHAPING_OUT, XNOR_1_6_N103_PULSESHAPING_OUT;
      NOR2_X1 XNOR_1_1_N103_PULSESHAPING (.ZN (XNOR_1_1_N103_PULSESHAPING_OUT), .A1 (N103_PWL), .A2 (GND));
      NOR2_X1 XNOR_1_2_N103_PULSESHAPING (.ZN (XNOR_1_2_N103_PULSESHAPING_OUT), .A1 (XNOR_1_1_N103_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_3_N103_PULSESHAPING (.ZN (XNOR_1_3_N103_PULSESHAPING_OUT), .A1 (XNOR_1_2_N103_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_4_N103_PULSESHAPING (.ZN (XNOR_1_4_N103_PULSESHAPING_OUT), .A1 (XNOR_1_3_N103_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_5_N103_PULSESHAPING (.ZN (XNOR_1_5_N103_PULSESHAPING_OUT), .A1 (XNOR_1_4_N103_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_6_N103_PULSESHAPING (.ZN (XNOR_1_6_N103_PULSESHAPING_OUT), .A1 (XNOR_1_5_N103_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_7_N103_PULSESHAPING (.ZN (N103), .A1 (XNOR_1_6_N103_PULSESHAPING_OUT), .A2 (GND));

      wire XNOR_1_1_N120_PULSESHAPING_OUT, XNOR_1_2_N120_PULSESHAPING_OUT, XNOR_1_3_N120_PULSESHAPING_OUT, XNOR_1_4_N120_PULSESHAPING_OUT, XNOR_1_5_N120_PULSESHAPING_OUT, XNOR_1_6_N120_PULSESHAPING_OUT;
      NOR2_X1 XNOR_1_1_N120_PULSESHAPING (.ZN (XNOR_1_1_N120_PULSESHAPING_OUT), .A1 (N120_PWL), .A2 (GND));
      NOR2_X1 XNOR_1_2_N120_PULSESHAPING (.ZN (XNOR_1_2_N120_PULSESHAPING_OUT), .A1 (XNOR_1_1_N120_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_3_N120_PULSESHAPING (.ZN (XNOR_1_3_N120_PULSESHAPING_OUT), .A1 (XNOR_1_2_N120_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_4_N120_PULSESHAPING (.ZN (XNOR_1_4_N120_PULSESHAPING_OUT), .A1 (XNOR_1_3_N120_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_5_N120_PULSESHAPING (.ZN (XNOR_1_5_N120_PULSESHAPING_OUT), .A1 (XNOR_1_4_N120_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_6_N120_PULSESHAPING (.ZN (XNOR_1_6_N120_PULSESHAPING_OUT), .A1 (XNOR_1_5_N120_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_7_N120_PULSESHAPING (.ZN (N120), .A1 (XNOR_1_6_N120_PULSESHAPING_OUT), .A2 (GND));

      wire XNOR_1_1_N137_PULSESHAPING_OUT, XNOR_1_2_N137_PULSESHAPING_OUT, XNOR_1_3_N137_PULSESHAPING_OUT, XNOR_1_4_N137_PULSESHAPING_OUT, XNOR_1_5_N137_PULSESHAPING_OUT, XNOR_1_6_N137_PULSESHAPING_OUT;
      NOR2_X1 XNOR_1_1_N137_PULSESHAPING (.ZN (XNOR_1_1_N137_PULSESHAPING_OUT), .A1 (N137_PWL), .A2 (GND));
      NOR2_X1 XNOR_1_2_N137_PULSESHAPING (.ZN (XNOR_1_2_N137_PULSESHAPING_OUT), .A1 (XNOR_1_1_N137_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_3_N137_PULSESHAPING (.ZN (XNOR_1_3_N137_PULSESHAPING_OUT), .A1 (XNOR_1_2_N137_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_4_N137_PULSESHAPING (.ZN (XNOR_1_4_N137_PULSESHAPING_OUT), .A1 (XNOR_1_3_N137_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_5_N137_PULSESHAPING (.ZN (XNOR_1_5_N137_PULSESHAPING_OUT), .A1 (XNOR_1_4_N137_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_6_N137_PULSESHAPING (.ZN (XNOR_1_6_N137_PULSESHAPING_OUT), .A1 (XNOR_1_5_N137_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_7_N137_PULSESHAPING (.ZN (N137), .A1 (XNOR_1_6_N137_PULSESHAPING_OUT), .A2 (GND));

      wire XNOR_1_1_N154_PULSESHAPING_OUT, XNOR_1_2_N154_PULSESHAPING_OUT, XNOR_1_3_N154_PULSESHAPING_OUT, XNOR_1_4_N154_PULSESHAPING_OUT, XNOR_1_5_N154_PULSESHAPING_OUT, XNOR_1_6_N154_PULSESHAPING_OUT;
      NOR2_X1 XNOR_1_1_N154_PULSESHAPING (.ZN (XNOR_1_1_N154_PULSESHAPING_OUT), .A1 (N154_PWL), .A2 (GND));
      NOR2_X1 XNOR_1_2_N154_PULSESHAPING (.ZN (XNOR_1_2_N154_PULSESHAPING_OUT), .A1 (XNOR_1_1_N154_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_3_N154_PULSESHAPING (.ZN (XNOR_1_3_N154_PULSESHAPING_OUT), .A1 (XNOR_1_2_N154_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_4_N154_PULSESHAPING (.ZN (XNOR_1_4_N154_PULSESHAPING_OUT), .A1 (XNOR_1_3_N154_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_5_N154_PULSESHAPING (.ZN (XNOR_1_5_N154_PULSESHAPING_OUT), .A1 (XNOR_1_4_N154_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_6_N154_PULSESHAPING (.ZN (XNOR_1_6_N154_PULSESHAPING_OUT), .A1 (XNOR_1_5_N154_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_7_N154_PULSESHAPING (.ZN (N154), .A1 (XNOR_1_6_N154_PULSESHAPING_OUT), .A2 (GND));

      wire XNOR_1_1_N171_PULSESHAPING_OUT, XNOR_1_2_N171_PULSESHAPING_OUT, XNOR_1_3_N171_PULSESHAPING_OUT, XNOR_1_4_N171_PULSESHAPING_OUT, XNOR_1_5_N171_PULSESHAPING_OUT, XNOR_1_6_N171_PULSESHAPING_OUT;
      NOR2_X1 XNOR_1_1_N171_PULSESHAPING (.ZN (XNOR_1_1_N171_PULSESHAPING_OUT), .A1 (N171_PWL), .A2 (GND));
      NOR2_X1 XNOR_1_2_N171_PULSESHAPING (.ZN (XNOR_1_2_N171_PULSESHAPING_OUT), .A1 (XNOR_1_1_N171_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_3_N171_PULSESHAPING (.ZN (XNOR_1_3_N171_PULSESHAPING_OUT), .A1 (XNOR_1_2_N171_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_4_N171_PULSESHAPING (.ZN (XNOR_1_4_N171_PULSESHAPING_OUT), .A1 (XNOR_1_3_N171_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_5_N171_PULSESHAPING (.ZN (XNOR_1_5_N171_PULSESHAPING_OUT), .A1 (XNOR_1_4_N171_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_6_N171_PULSESHAPING (.ZN (XNOR_1_6_N171_PULSESHAPING_OUT), .A1 (XNOR_1_5_N171_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_7_N171_PULSESHAPING (.ZN (N171), .A1 (XNOR_1_6_N171_PULSESHAPING_OUT), .A2 (GND));

      wire XNOR_1_1_N188_PULSESHAPING_OUT, XNOR_1_2_N188_PULSESHAPING_OUT, XNOR_1_3_N188_PULSESHAPING_OUT, XNOR_1_4_N188_PULSESHAPING_OUT, XNOR_1_5_N188_PULSESHAPING_OUT, XNOR_1_6_N188_PULSESHAPING_OUT;
      NOR2_X1 XNOR_1_1_N188_PULSESHAPING (.ZN (XNOR_1_1_N188_PULSESHAPING_OUT), .A1 (N188_PWL), .A2 (GND));
      NOR2_X1 XNOR_1_2_N188_PULSESHAPING (.ZN (XNOR_1_2_N188_PULSESHAPING_OUT), .A1 (XNOR_1_1_N188_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_3_N188_PULSESHAPING (.ZN (XNOR_1_3_N188_PULSESHAPING_OUT), .A1 (XNOR_1_2_N188_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_4_N188_PULSESHAPING (.ZN (XNOR_1_4_N188_PULSESHAPING_OUT), .A1 (XNOR_1_3_N188_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_5_N188_PULSESHAPING (.ZN (XNOR_1_5_N188_PULSESHAPING_OUT), .A1 (XNOR_1_4_N188_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_6_N188_PULSESHAPING (.ZN (XNOR_1_6_N188_PULSESHAPING_OUT), .A1 (XNOR_1_5_N188_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_7_N188_PULSESHAPING (.ZN (N188), .A1 (XNOR_1_6_N188_PULSESHAPING_OUT), .A2 (GND));

      wire XNOR_1_1_N205_PULSESHAPING_OUT, XNOR_1_2_N205_PULSESHAPING_OUT, XNOR_1_3_N205_PULSESHAPING_OUT, XNOR_1_4_N205_PULSESHAPING_OUT, XNOR_1_5_N205_PULSESHAPING_OUT, XNOR_1_6_N205_PULSESHAPING_OUT;
      NOR2_X1 XNOR_1_1_N205_PULSESHAPING (.ZN (XNOR_1_1_N205_PULSESHAPING_OUT), .A1 (N205_PWL), .A2 (GND));
      NOR2_X1 XNOR_1_2_N205_PULSESHAPING (.ZN (XNOR_1_2_N205_PULSESHAPING_OUT), .A1 (XNOR_1_1_N205_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_3_N205_PULSESHAPING (.ZN (XNOR_1_3_N205_PULSESHAPING_OUT), .A1 (XNOR_1_2_N205_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_4_N205_PULSESHAPING (.ZN (XNOR_1_4_N205_PULSESHAPING_OUT), .A1 (XNOR_1_3_N205_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_5_N205_PULSESHAPING (.ZN (XNOR_1_5_N205_PULSESHAPING_OUT), .A1 (XNOR_1_4_N205_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_6_N205_PULSESHAPING (.ZN (XNOR_1_6_N205_PULSESHAPING_OUT), .A1 (XNOR_1_5_N205_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_7_N205_PULSESHAPING (.ZN (N205), .A1 (XNOR_1_6_N205_PULSESHAPING_OUT), .A2 (GND));

      wire XNOR_1_1_N222_PULSESHAPING_OUT, XNOR_1_2_N222_PULSESHAPING_OUT, XNOR_1_3_N222_PULSESHAPING_OUT, XNOR_1_4_N222_PULSESHAPING_OUT, XNOR_1_5_N222_PULSESHAPING_OUT, XNOR_1_6_N222_PULSESHAPING_OUT;
      NOR2_X1 XNOR_1_1_N222_PULSESHAPING (.ZN (XNOR_1_1_N222_PULSESHAPING_OUT), .A1 (N222_PWL), .A2 (GND));
      NOR2_X1 XNOR_1_2_N222_PULSESHAPING (.ZN (XNOR_1_2_N222_PULSESHAPING_OUT), .A1 (XNOR_1_1_N222_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_3_N222_PULSESHAPING (.ZN (XNOR_1_3_N222_PULSESHAPING_OUT), .A1 (XNOR_1_2_N222_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_4_N222_PULSESHAPING (.ZN (XNOR_1_4_N222_PULSESHAPING_OUT), .A1 (XNOR_1_3_N222_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_5_N222_PULSESHAPING (.ZN (XNOR_1_5_N222_PULSESHAPING_OUT), .A1 (XNOR_1_4_N222_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_6_N222_PULSESHAPING (.ZN (XNOR_1_6_N222_PULSESHAPING_OUT), .A1 (XNOR_1_5_N222_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_7_N222_PULSESHAPING (.ZN (N222), .A1 (XNOR_1_6_N222_PULSESHAPING_OUT), .A2 (GND));

      wire XNOR_1_1_N239_PULSESHAPING_OUT, XNOR_1_2_N239_PULSESHAPING_OUT, XNOR_1_3_N239_PULSESHAPING_OUT, XNOR_1_4_N239_PULSESHAPING_OUT, XNOR_1_5_N239_PULSESHAPING_OUT, XNOR_1_6_N239_PULSESHAPING_OUT;
      NOR2_X1 XNOR_1_1_N239_PULSESHAPING (.ZN (XNOR_1_1_N239_PULSESHAPING_OUT), .A1 (N239_PWL), .A2 (GND));
      NOR2_X1 XNOR_1_2_N239_PULSESHAPING (.ZN (XNOR_1_2_N239_PULSESHAPING_OUT), .A1 (XNOR_1_1_N239_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_3_N239_PULSESHAPING (.ZN (XNOR_1_3_N239_PULSESHAPING_OUT), .A1 (XNOR_1_2_N239_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_4_N239_PULSESHAPING (.ZN (XNOR_1_4_N239_PULSESHAPING_OUT), .A1 (XNOR_1_3_N239_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_5_N239_PULSESHAPING (.ZN (XNOR_1_5_N239_PULSESHAPING_OUT), .A1 (XNOR_1_4_N239_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_6_N239_PULSESHAPING (.ZN (XNOR_1_6_N239_PULSESHAPING_OUT), .A1 (XNOR_1_5_N239_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_7_N239_PULSESHAPING (.ZN (N239), .A1 (XNOR_1_6_N239_PULSESHAPING_OUT), .A2 (GND));

      wire XNOR_1_1_N256_PULSESHAPING_OUT, XNOR_1_2_N256_PULSESHAPING_OUT, XNOR_1_3_N256_PULSESHAPING_OUT, XNOR_1_4_N256_PULSESHAPING_OUT, XNOR_1_5_N256_PULSESHAPING_OUT, XNOR_1_6_N256_PULSESHAPING_OUT;
      NOR2_X1 XNOR_1_1_N256_PULSESHAPING (.ZN (XNOR_1_1_N256_PULSESHAPING_OUT), .A1 (N256_PWL), .A2 (GND));
      NOR2_X1 XNOR_1_2_N256_PULSESHAPING (.ZN (XNOR_1_2_N256_PULSESHAPING_OUT), .A1 (XNOR_1_1_N256_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_3_N256_PULSESHAPING (.ZN (XNOR_1_3_N256_PULSESHAPING_OUT), .A1 (XNOR_1_2_N256_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_4_N256_PULSESHAPING (.ZN (XNOR_1_4_N256_PULSESHAPING_OUT), .A1 (XNOR_1_3_N256_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_5_N256_PULSESHAPING (.ZN (XNOR_1_5_N256_PULSESHAPING_OUT), .A1 (XNOR_1_4_N256_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_6_N256_PULSESHAPING (.ZN (XNOR_1_6_N256_PULSESHAPING_OUT), .A1 (XNOR_1_5_N256_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_7_N256_PULSESHAPING (.ZN (N256), .A1 (XNOR_1_6_N256_PULSESHAPING_OUT), .A2 (GND));

      wire XNOR_1_1_N273_PULSESHAPING_OUT, XNOR_1_2_N273_PULSESHAPING_OUT, XNOR_1_3_N273_PULSESHAPING_OUT, XNOR_1_4_N273_PULSESHAPING_OUT, XNOR_1_5_N273_PULSESHAPING_OUT, XNOR_1_6_N273_PULSESHAPING_OUT;
      NOR2_X1 XNOR_1_1_N273_PULSESHAPING (.ZN (XNOR_1_1_N273_PULSESHAPING_OUT), .A1 (N273_PWL), .A2 (GND));
      NOR2_X1 XNOR_1_2_N273_PULSESHAPING (.ZN (XNOR_1_2_N273_PULSESHAPING_OUT), .A1 (XNOR_1_1_N273_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_3_N273_PULSESHAPING (.ZN (XNOR_1_3_N273_PULSESHAPING_OUT), .A1 (XNOR_1_2_N273_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_4_N273_PULSESHAPING (.ZN (XNOR_1_4_N273_PULSESHAPING_OUT), .A1 (XNOR_1_3_N273_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_5_N273_PULSESHAPING (.ZN (XNOR_1_5_N273_PULSESHAPING_OUT), .A1 (XNOR_1_4_N273_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_6_N273_PULSESHAPING (.ZN (XNOR_1_6_N273_PULSESHAPING_OUT), .A1 (XNOR_1_5_N273_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_7_N273_PULSESHAPING (.ZN (N273), .A1 (XNOR_1_6_N273_PULSESHAPING_OUT), .A2 (GND));

      wire XNOR_1_1_N290_PULSESHAPING_OUT, XNOR_1_2_N290_PULSESHAPING_OUT, XNOR_1_3_N290_PULSESHAPING_OUT, XNOR_1_4_N290_PULSESHAPING_OUT, XNOR_1_5_N290_PULSESHAPING_OUT, XNOR_1_6_N290_PULSESHAPING_OUT;
      NOR2_X1 XNOR_1_1_N290_PULSESHAPING (.ZN (XNOR_1_1_N290_PULSESHAPING_OUT), .A1 (N290_PWL), .A2 (GND));
      NOR2_X1 XNOR_1_2_N290_PULSESHAPING (.ZN (XNOR_1_2_N290_PULSESHAPING_OUT), .A1 (XNOR_1_1_N290_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_3_N290_PULSESHAPING (.ZN (XNOR_1_3_N290_PULSESHAPING_OUT), .A1 (XNOR_1_2_N290_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_4_N290_PULSESHAPING (.ZN (XNOR_1_4_N290_PULSESHAPING_OUT), .A1 (XNOR_1_3_N290_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_5_N290_PULSESHAPING (.ZN (XNOR_1_5_N290_PULSESHAPING_OUT), .A1 (XNOR_1_4_N290_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_6_N290_PULSESHAPING (.ZN (XNOR_1_6_N290_PULSESHAPING_OUT), .A1 (XNOR_1_5_N290_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_7_N290_PULSESHAPING (.ZN (N290), .A1 (XNOR_1_6_N290_PULSESHAPING_OUT), .A2 (GND));

      wire XNOR_1_1_N307_PULSESHAPING_OUT, XNOR_1_2_N307_PULSESHAPING_OUT, XNOR_1_3_N307_PULSESHAPING_OUT, XNOR_1_4_N307_PULSESHAPING_OUT, XNOR_1_5_N307_PULSESHAPING_OUT, XNOR_1_6_N307_PULSESHAPING_OUT;
      NOR2_X1 XNOR_1_1_N307_PULSESHAPING (.ZN (XNOR_1_1_N307_PULSESHAPING_OUT), .A1 (N307_PWL), .A2 (GND));
      NOR2_X1 XNOR_1_2_N307_PULSESHAPING (.ZN (XNOR_1_2_N307_PULSESHAPING_OUT), .A1 (XNOR_1_1_N307_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_3_N307_PULSESHAPING (.ZN (XNOR_1_3_N307_PULSESHAPING_OUT), .A1 (XNOR_1_2_N307_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_4_N307_PULSESHAPING (.ZN (XNOR_1_4_N307_PULSESHAPING_OUT), .A1 (XNOR_1_3_N307_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_5_N307_PULSESHAPING (.ZN (XNOR_1_5_N307_PULSESHAPING_OUT), .A1 (XNOR_1_4_N307_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_6_N307_PULSESHAPING (.ZN (XNOR_1_6_N307_PULSESHAPING_OUT), .A1 (XNOR_1_5_N307_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_7_N307_PULSESHAPING (.ZN (N307), .A1 (XNOR_1_6_N307_PULSESHAPING_OUT), .A2 (GND));

      wire XNOR_1_1_N324_PULSESHAPING_OUT, XNOR_1_2_N324_PULSESHAPING_OUT, XNOR_1_3_N324_PULSESHAPING_OUT, XNOR_1_4_N324_PULSESHAPING_OUT, XNOR_1_5_N324_PULSESHAPING_OUT, XNOR_1_6_N324_PULSESHAPING_OUT;
      NOR2_X1 XNOR_1_1_N324_PULSESHAPING (.ZN (XNOR_1_1_N324_PULSESHAPING_OUT), .A1 (N324_PWL), .A2 (GND));
      NOR2_X1 XNOR_1_2_N324_PULSESHAPING (.ZN (XNOR_1_2_N324_PULSESHAPING_OUT), .A1 (XNOR_1_1_N324_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_3_N324_PULSESHAPING (.ZN (XNOR_1_3_N324_PULSESHAPING_OUT), .A1 (XNOR_1_2_N324_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_4_N324_PULSESHAPING (.ZN (XNOR_1_4_N324_PULSESHAPING_OUT), .A1 (XNOR_1_3_N324_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_5_N324_PULSESHAPING (.ZN (XNOR_1_5_N324_PULSESHAPING_OUT), .A1 (XNOR_1_4_N324_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_6_N324_PULSESHAPING (.ZN (XNOR_1_6_N324_PULSESHAPING_OUT), .A1 (XNOR_1_5_N324_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_7_N324_PULSESHAPING (.ZN (N324), .A1 (XNOR_1_6_N324_PULSESHAPING_OUT), .A2 (GND));

      wire XNOR_1_1_N341_PULSESHAPING_OUT, XNOR_1_2_N341_PULSESHAPING_OUT, XNOR_1_3_N341_PULSESHAPING_OUT, XNOR_1_4_N341_PULSESHAPING_OUT, XNOR_1_5_N341_PULSESHAPING_OUT, XNOR_1_6_N341_PULSESHAPING_OUT;
      NOR2_X1 XNOR_1_1_N341_PULSESHAPING (.ZN (XNOR_1_1_N341_PULSESHAPING_OUT), .A1 (N341_PWL), .A2 (GND));
      NOR2_X1 XNOR_1_2_N341_PULSESHAPING (.ZN (XNOR_1_2_N341_PULSESHAPING_OUT), .A1 (XNOR_1_1_N341_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_3_N341_PULSESHAPING (.ZN (XNOR_1_3_N341_PULSESHAPING_OUT), .A1 (XNOR_1_2_N341_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_4_N341_PULSESHAPING (.ZN (XNOR_1_4_N341_PULSESHAPING_OUT), .A1 (XNOR_1_3_N341_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_5_N341_PULSESHAPING (.ZN (XNOR_1_5_N341_PULSESHAPING_OUT), .A1 (XNOR_1_4_N341_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_6_N341_PULSESHAPING (.ZN (XNOR_1_6_N341_PULSESHAPING_OUT), .A1 (XNOR_1_5_N341_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_7_N341_PULSESHAPING (.ZN (N341), .A1 (XNOR_1_6_N341_PULSESHAPING_OUT), .A2 (GND));

      wire XNOR_1_1_N358_PULSESHAPING_OUT, XNOR_1_2_N358_PULSESHAPING_OUT, XNOR_1_3_N358_PULSESHAPING_OUT, XNOR_1_4_N358_PULSESHAPING_OUT, XNOR_1_5_N358_PULSESHAPING_OUT, XNOR_1_6_N358_PULSESHAPING_OUT;
      NOR2_X1 XNOR_1_1_N358_PULSESHAPING (.ZN (XNOR_1_1_N358_PULSESHAPING_OUT), .A1 (N358_PWL), .A2 (GND));
      NOR2_X1 XNOR_1_2_N358_PULSESHAPING (.ZN (XNOR_1_2_N358_PULSESHAPING_OUT), .A1 (XNOR_1_1_N358_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_3_N358_PULSESHAPING (.ZN (XNOR_1_3_N358_PULSESHAPING_OUT), .A1 (XNOR_1_2_N358_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_4_N358_PULSESHAPING (.ZN (XNOR_1_4_N358_PULSESHAPING_OUT), .A1 (XNOR_1_3_N358_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_5_N358_PULSESHAPING (.ZN (XNOR_1_5_N358_PULSESHAPING_OUT), .A1 (XNOR_1_4_N358_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_6_N358_PULSESHAPING (.ZN (XNOR_1_6_N358_PULSESHAPING_OUT), .A1 (XNOR_1_5_N358_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_7_N358_PULSESHAPING (.ZN (N358), .A1 (XNOR_1_6_N358_PULSESHAPING_OUT), .A2 (GND));

      wire XNOR_1_1_N375_PULSESHAPING_OUT, XNOR_1_2_N375_PULSESHAPING_OUT, XNOR_1_3_N375_PULSESHAPING_OUT, XNOR_1_4_N375_PULSESHAPING_OUT, XNOR_1_5_N375_PULSESHAPING_OUT, XNOR_1_6_N375_PULSESHAPING_OUT;
      NOR2_X1 XNOR_1_1_N375_PULSESHAPING (.ZN (XNOR_1_1_N375_PULSESHAPING_OUT), .A1 (N375_PWL), .A2 (GND));
      NOR2_X1 XNOR_1_2_N375_PULSESHAPING (.ZN (XNOR_1_2_N375_PULSESHAPING_OUT), .A1 (XNOR_1_1_N375_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_3_N375_PULSESHAPING (.ZN (XNOR_1_3_N375_PULSESHAPING_OUT), .A1 (XNOR_1_2_N375_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_4_N375_PULSESHAPING (.ZN (XNOR_1_4_N375_PULSESHAPING_OUT), .A1 (XNOR_1_3_N375_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_5_N375_PULSESHAPING (.ZN (XNOR_1_5_N375_PULSESHAPING_OUT), .A1 (XNOR_1_4_N375_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_6_N375_PULSESHAPING (.ZN (XNOR_1_6_N375_PULSESHAPING_OUT), .A1 (XNOR_1_5_N375_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_7_N375_PULSESHAPING (.ZN (N375), .A1 (XNOR_1_6_N375_PULSESHAPING_OUT), .A2 (GND));

      wire XNOR_1_1_N392_PULSESHAPING_OUT, XNOR_1_2_N392_PULSESHAPING_OUT, XNOR_1_3_N392_PULSESHAPING_OUT, XNOR_1_4_N392_PULSESHAPING_OUT, XNOR_1_5_N392_PULSESHAPING_OUT, XNOR_1_6_N392_PULSESHAPING_OUT;
      NOR2_X1 XNOR_1_1_N392_PULSESHAPING (.ZN (XNOR_1_1_N392_PULSESHAPING_OUT), .A1 (N392_PWL), .A2 (GND));
      NOR2_X1 XNOR_1_2_N392_PULSESHAPING (.ZN (XNOR_1_2_N392_PULSESHAPING_OUT), .A1 (XNOR_1_1_N392_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_3_N392_PULSESHAPING (.ZN (XNOR_1_3_N392_PULSESHAPING_OUT), .A1 (XNOR_1_2_N392_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_4_N392_PULSESHAPING (.ZN (XNOR_1_4_N392_PULSESHAPING_OUT), .A1 (XNOR_1_3_N392_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_5_N392_PULSESHAPING (.ZN (XNOR_1_5_N392_PULSESHAPING_OUT), .A1 (XNOR_1_4_N392_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_6_N392_PULSESHAPING (.ZN (XNOR_1_6_N392_PULSESHAPING_OUT), .A1 (XNOR_1_5_N392_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_7_N392_PULSESHAPING (.ZN (N392), .A1 (XNOR_1_6_N392_PULSESHAPING_OUT), .A2 (GND));

      wire XNOR_1_1_N409_PULSESHAPING_OUT, XNOR_1_2_N409_PULSESHAPING_OUT, XNOR_1_3_N409_PULSESHAPING_OUT, XNOR_1_4_N409_PULSESHAPING_OUT, XNOR_1_5_N409_PULSESHAPING_OUT, XNOR_1_6_N409_PULSESHAPING_OUT;
      NOR2_X1 XNOR_1_1_N409_PULSESHAPING (.ZN (XNOR_1_1_N409_PULSESHAPING_OUT), .A1 (N409_PWL), .A2 (GND));
      NOR2_X1 XNOR_1_2_N409_PULSESHAPING (.ZN (XNOR_1_2_N409_PULSESHAPING_OUT), .A1 (XNOR_1_1_N409_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_3_N409_PULSESHAPING (.ZN (XNOR_1_3_N409_PULSESHAPING_OUT), .A1 (XNOR_1_2_N409_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_4_N409_PULSESHAPING (.ZN (XNOR_1_4_N409_PULSESHAPING_OUT), .A1 (XNOR_1_3_N409_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_5_N409_PULSESHAPING (.ZN (XNOR_1_5_N409_PULSESHAPING_OUT), .A1 (XNOR_1_4_N409_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_6_N409_PULSESHAPING (.ZN (XNOR_1_6_N409_PULSESHAPING_OUT), .A1 (XNOR_1_5_N409_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_7_N409_PULSESHAPING (.ZN (N409), .A1 (XNOR_1_6_N409_PULSESHAPING_OUT), .A2 (GND));

      wire XNOR_1_1_N426_PULSESHAPING_OUT, XNOR_1_2_N426_PULSESHAPING_OUT, XNOR_1_3_N426_PULSESHAPING_OUT, XNOR_1_4_N426_PULSESHAPING_OUT, XNOR_1_5_N426_PULSESHAPING_OUT, XNOR_1_6_N426_PULSESHAPING_OUT;
      NOR2_X1 XNOR_1_1_N426_PULSESHAPING (.ZN (XNOR_1_1_N426_PULSESHAPING_OUT), .A1 (N426_PWL), .A2 (GND));
      NOR2_X1 XNOR_1_2_N426_PULSESHAPING (.ZN (XNOR_1_2_N426_PULSESHAPING_OUT), .A1 (XNOR_1_1_N426_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_3_N426_PULSESHAPING (.ZN (XNOR_1_3_N426_PULSESHAPING_OUT), .A1 (XNOR_1_2_N426_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_4_N426_PULSESHAPING (.ZN (XNOR_1_4_N426_PULSESHAPING_OUT), .A1 (XNOR_1_3_N426_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_5_N426_PULSESHAPING (.ZN (XNOR_1_5_N426_PULSESHAPING_OUT), .A1 (XNOR_1_4_N426_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_6_N426_PULSESHAPING (.ZN (XNOR_1_6_N426_PULSESHAPING_OUT), .A1 (XNOR_1_5_N426_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_7_N426_PULSESHAPING (.ZN (N426), .A1 (XNOR_1_6_N426_PULSESHAPING_OUT), .A2 (GND));

      wire XNOR_1_1_N443_PULSESHAPING_OUT, XNOR_1_2_N443_PULSESHAPING_OUT, XNOR_1_3_N443_PULSESHAPING_OUT, XNOR_1_4_N443_PULSESHAPING_OUT, XNOR_1_5_N443_PULSESHAPING_OUT, XNOR_1_6_N443_PULSESHAPING_OUT;
      NOR2_X1 XNOR_1_1_N443_PULSESHAPING (.ZN (XNOR_1_1_N443_PULSESHAPING_OUT), .A1 (N443_PWL), .A2 (GND));
      NOR2_X1 XNOR_1_2_N443_PULSESHAPING (.ZN (XNOR_1_2_N443_PULSESHAPING_OUT), .A1 (XNOR_1_1_N443_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_3_N443_PULSESHAPING (.ZN (XNOR_1_3_N443_PULSESHAPING_OUT), .A1 (XNOR_1_2_N443_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_4_N443_PULSESHAPING (.ZN (XNOR_1_4_N443_PULSESHAPING_OUT), .A1 (XNOR_1_3_N443_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_5_N443_PULSESHAPING (.ZN (XNOR_1_5_N443_PULSESHAPING_OUT), .A1 (XNOR_1_4_N443_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_6_N443_PULSESHAPING (.ZN (XNOR_1_6_N443_PULSESHAPING_OUT), .A1 (XNOR_1_5_N443_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_7_N443_PULSESHAPING (.ZN (N443), .A1 (XNOR_1_6_N443_PULSESHAPING_OUT), .A2 (GND));

      wire XNOR_1_1_N460_PULSESHAPING_OUT, XNOR_1_2_N460_PULSESHAPING_OUT, XNOR_1_3_N460_PULSESHAPING_OUT, XNOR_1_4_N460_PULSESHAPING_OUT, XNOR_1_5_N460_PULSESHAPING_OUT, XNOR_1_6_N460_PULSESHAPING_OUT;
      NOR2_X1 XNOR_1_1_N460_PULSESHAPING (.ZN (XNOR_1_1_N460_PULSESHAPING_OUT), .A1 (N460_PWL), .A2 (GND));
      NOR2_X1 XNOR_1_2_N460_PULSESHAPING (.ZN (XNOR_1_2_N460_PULSESHAPING_OUT), .A1 (XNOR_1_1_N460_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_3_N460_PULSESHAPING (.ZN (XNOR_1_3_N460_PULSESHAPING_OUT), .A1 (XNOR_1_2_N460_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_4_N460_PULSESHAPING (.ZN (XNOR_1_4_N460_PULSESHAPING_OUT), .A1 (XNOR_1_3_N460_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_5_N460_PULSESHAPING (.ZN (XNOR_1_5_N460_PULSESHAPING_OUT), .A1 (XNOR_1_4_N460_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_6_N460_PULSESHAPING (.ZN (XNOR_1_6_N460_PULSESHAPING_OUT), .A1 (XNOR_1_5_N460_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_7_N460_PULSESHAPING (.ZN (N460), .A1 (XNOR_1_6_N460_PULSESHAPING_OUT), .A2 (GND));

      wire XNOR_1_1_N477_PULSESHAPING_OUT, XNOR_1_2_N477_PULSESHAPING_OUT, XNOR_1_3_N477_PULSESHAPING_OUT, XNOR_1_4_N477_PULSESHAPING_OUT, XNOR_1_5_N477_PULSESHAPING_OUT, XNOR_1_6_N477_PULSESHAPING_OUT;
      NOR2_X1 XNOR_1_1_N477_PULSESHAPING (.ZN (XNOR_1_1_N477_PULSESHAPING_OUT), .A1 (N477_PWL), .A2 (GND));
      NOR2_X1 XNOR_1_2_N477_PULSESHAPING (.ZN (XNOR_1_2_N477_PULSESHAPING_OUT), .A1 (XNOR_1_1_N477_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_3_N477_PULSESHAPING (.ZN (XNOR_1_3_N477_PULSESHAPING_OUT), .A1 (XNOR_1_2_N477_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_4_N477_PULSESHAPING (.ZN (XNOR_1_4_N477_PULSESHAPING_OUT), .A1 (XNOR_1_3_N477_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_5_N477_PULSESHAPING (.ZN (XNOR_1_5_N477_PULSESHAPING_OUT), .A1 (XNOR_1_4_N477_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_6_N477_PULSESHAPING (.ZN (XNOR_1_6_N477_PULSESHAPING_OUT), .A1 (XNOR_1_5_N477_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_7_N477_PULSESHAPING (.ZN (N477), .A1 (XNOR_1_6_N477_PULSESHAPING_OUT), .A2 (GND));

      wire XNOR_1_1_N494_PULSESHAPING_OUT, XNOR_1_2_N494_PULSESHAPING_OUT, XNOR_1_3_N494_PULSESHAPING_OUT, XNOR_1_4_N494_PULSESHAPING_OUT, XNOR_1_5_N494_PULSESHAPING_OUT, XNOR_1_6_N494_PULSESHAPING_OUT;
      NOR2_X1 XNOR_1_1_N494_PULSESHAPING (.ZN (XNOR_1_1_N494_PULSESHAPING_OUT), .A1 (N494_PWL), .A2 (GND));
      NOR2_X1 XNOR_1_2_N494_PULSESHAPING (.ZN (XNOR_1_2_N494_PULSESHAPING_OUT), .A1 (XNOR_1_1_N494_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_3_N494_PULSESHAPING (.ZN (XNOR_1_3_N494_PULSESHAPING_OUT), .A1 (XNOR_1_2_N494_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_4_N494_PULSESHAPING (.ZN (XNOR_1_4_N494_PULSESHAPING_OUT), .A1 (XNOR_1_3_N494_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_5_N494_PULSESHAPING (.ZN (XNOR_1_5_N494_PULSESHAPING_OUT), .A1 (XNOR_1_4_N494_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_6_N494_PULSESHAPING (.ZN (XNOR_1_6_N494_PULSESHAPING_OUT), .A1 (XNOR_1_5_N494_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_7_N494_PULSESHAPING (.ZN (N494), .A1 (XNOR_1_6_N494_PULSESHAPING_OUT), .A2 (GND));

      wire XNOR_1_1_N511_PULSESHAPING_OUT, XNOR_1_2_N511_PULSESHAPING_OUT, XNOR_1_3_N511_PULSESHAPING_OUT, XNOR_1_4_N511_PULSESHAPING_OUT, XNOR_1_5_N511_PULSESHAPING_OUT, XNOR_1_6_N511_PULSESHAPING_OUT;
      NOR2_X1 XNOR_1_1_N511_PULSESHAPING (.ZN (XNOR_1_1_N511_PULSESHAPING_OUT), .A1 (N511_PWL), .A2 (GND));
      NOR2_X1 XNOR_1_2_N511_PULSESHAPING (.ZN (XNOR_1_2_N511_PULSESHAPING_OUT), .A1 (XNOR_1_1_N511_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_3_N511_PULSESHAPING (.ZN (XNOR_1_3_N511_PULSESHAPING_OUT), .A1 (XNOR_1_2_N511_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_4_N511_PULSESHAPING (.ZN (XNOR_1_4_N511_PULSESHAPING_OUT), .A1 (XNOR_1_3_N511_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_5_N511_PULSESHAPING (.ZN (XNOR_1_5_N511_PULSESHAPING_OUT), .A1 (XNOR_1_4_N511_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_6_N511_PULSESHAPING (.ZN (XNOR_1_6_N511_PULSESHAPING_OUT), .A1 (XNOR_1_5_N511_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_7_N511_PULSESHAPING (.ZN (N511), .A1 (XNOR_1_6_N511_PULSESHAPING_OUT), .A2 (GND));

      wire XNOR_1_1_N528_PULSESHAPING_OUT, XNOR_1_2_N528_PULSESHAPING_OUT, XNOR_1_3_N528_PULSESHAPING_OUT, XNOR_1_4_N528_PULSESHAPING_OUT, XNOR_1_5_N528_PULSESHAPING_OUT, XNOR_1_6_N528_PULSESHAPING_OUT;
      NOR2_X1 XNOR_1_1_N528_PULSESHAPING (.ZN (XNOR_1_1_N528_PULSESHAPING_OUT), .A1 (N528_PWL), .A2 (GND));
      NOR2_X1 XNOR_1_2_N528_PULSESHAPING (.ZN (XNOR_1_2_N528_PULSESHAPING_OUT), .A1 (XNOR_1_1_N528_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_3_N528_PULSESHAPING (.ZN (XNOR_1_3_N528_PULSESHAPING_OUT), .A1 (XNOR_1_2_N528_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_4_N528_PULSESHAPING (.ZN (XNOR_1_4_N528_PULSESHAPING_OUT), .A1 (XNOR_1_3_N528_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_5_N528_PULSESHAPING (.ZN (XNOR_1_5_N528_PULSESHAPING_OUT), .A1 (XNOR_1_4_N528_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_6_N528_PULSESHAPING (.ZN (XNOR_1_6_N528_PULSESHAPING_OUT), .A1 (XNOR_1_5_N528_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_7_N528_PULSESHAPING (.ZN (N528), .A1 (XNOR_1_6_N528_PULSESHAPING_OUT), .A2 (GND));



      wire XNOR_1_1_AND2_NUM1_OUT, XNOR_1_2_AND2_NUM1_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM1 (.ZN (XNOR_1_1_AND2_NUM1_OUT), .A1 (N1), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM1 (.ZN (XNOR_1_2_AND2_NUM1_OUT), .A1 (GND), .A2 (N273));
      NOR2_X1 XNOR_1_3_AND2_NUM1 (.ZN (N545), .A1 (XNOR_1_1_AND2_NUM1_OUT), .A2 (XNOR_1_2_AND2_NUM1_OUT));
      wire XNOR_1_1_AND2_NUM2_OUT, XNOR_1_2_AND2_NUM2_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM2 (.ZN (XNOR_1_1_AND2_NUM2_OUT), .A1 (N1), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM2 (.ZN (XNOR_1_2_AND2_NUM2_OUT), .A1 (GND), .A2 (N290));
      NOR2_X1 XNOR_1_3_AND2_NUM2 (.ZN (N546), .A1 (XNOR_1_1_AND2_NUM2_OUT), .A2 (XNOR_1_2_AND2_NUM2_OUT));
      wire XNOR_1_1_AND2_NUM3_OUT, XNOR_1_2_AND2_NUM3_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM3 (.ZN (XNOR_1_1_AND2_NUM3_OUT), .A1 (N1), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM3 (.ZN (XNOR_1_2_AND2_NUM3_OUT), .A1 (GND), .A2 (N307));
      NOR2_X1 XNOR_1_3_AND2_NUM3 (.ZN (N549), .A1 (XNOR_1_1_AND2_NUM3_OUT), .A2 (XNOR_1_2_AND2_NUM3_OUT));
      wire XNOR_1_1_AND2_NUM4_OUT, XNOR_1_2_AND2_NUM4_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM4 (.ZN (XNOR_1_1_AND2_NUM4_OUT), .A1 (N1), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM4 (.ZN (XNOR_1_2_AND2_NUM4_OUT), .A1 (GND), .A2 (N324));
      NOR2_X1 XNOR_1_3_AND2_NUM4 (.ZN (N552), .A1 (XNOR_1_1_AND2_NUM4_OUT), .A2 (XNOR_1_2_AND2_NUM4_OUT));
      wire XNOR_1_1_AND2_NUM5_OUT, XNOR_1_2_AND2_NUM5_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM5 (.ZN (XNOR_1_1_AND2_NUM5_OUT), .A1 (N1), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM5 (.ZN (XNOR_1_2_AND2_NUM5_OUT), .A1 (GND), .A2 (N341));
      NOR2_X1 XNOR_1_3_AND2_NUM5 (.ZN (N555), .A1 (XNOR_1_1_AND2_NUM5_OUT), .A2 (XNOR_1_2_AND2_NUM5_OUT));
      wire XNOR_1_1_AND2_NUM6_OUT, XNOR_1_2_AND2_NUM6_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM6 (.ZN (XNOR_1_1_AND2_NUM6_OUT), .A1 (N1), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM6 (.ZN (XNOR_1_2_AND2_NUM6_OUT), .A1 (GND), .A2 (N358));
      NOR2_X1 XNOR_1_3_AND2_NUM6 (.ZN (N558), .A1 (XNOR_1_1_AND2_NUM6_OUT), .A2 (XNOR_1_2_AND2_NUM6_OUT));
      wire XNOR_1_1_AND2_NUM7_OUT, XNOR_1_2_AND2_NUM7_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM7 (.ZN (XNOR_1_1_AND2_NUM7_OUT), .A1 (N1), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM7 (.ZN (XNOR_1_2_AND2_NUM7_OUT), .A1 (GND), .A2 (N375));
      NOR2_X1 XNOR_1_3_AND2_NUM7 (.ZN (N561), .A1 (XNOR_1_1_AND2_NUM7_OUT), .A2 (XNOR_1_2_AND2_NUM7_OUT));
      wire XNOR_1_1_AND2_NUM8_OUT, XNOR_1_2_AND2_NUM8_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM8 (.ZN (XNOR_1_1_AND2_NUM8_OUT), .A1 (N1), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM8 (.ZN (XNOR_1_2_AND2_NUM8_OUT), .A1 (GND), .A2 (N392));
      NOR2_X1 XNOR_1_3_AND2_NUM8 (.ZN (N564), .A1 (XNOR_1_1_AND2_NUM8_OUT), .A2 (XNOR_1_2_AND2_NUM8_OUT));
      wire XNOR_1_1_AND2_NUM9_OUT, XNOR_1_2_AND2_NUM9_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM9 (.ZN (XNOR_1_1_AND2_NUM9_OUT), .A1 (N1), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM9 (.ZN (XNOR_1_2_AND2_NUM9_OUT), .A1 (GND), .A2 (N409));
      NOR2_X1 XNOR_1_3_AND2_NUM9 (.ZN (N567), .A1 (XNOR_1_1_AND2_NUM9_OUT), .A2 (XNOR_1_2_AND2_NUM9_OUT));
      wire XNOR_1_1_AND2_NUM10_OUT, XNOR_1_2_AND2_NUM10_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM10 (.ZN (XNOR_1_1_AND2_NUM10_OUT), .A1 (N1), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM10 (.ZN (XNOR_1_2_AND2_NUM10_OUT), .A1 (GND), .A2 (N426));
      NOR2_X1 XNOR_1_3_AND2_NUM10 (.ZN (N570), .A1 (XNOR_1_1_AND2_NUM10_OUT), .A2 (XNOR_1_2_AND2_NUM10_OUT));
      wire XNOR_1_1_AND2_NUM11_OUT, XNOR_1_2_AND2_NUM11_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM11 (.ZN (XNOR_1_1_AND2_NUM11_OUT), .A1 (N1), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM11 (.ZN (XNOR_1_2_AND2_NUM11_OUT), .A1 (GND), .A2 (N443));
      NOR2_X1 XNOR_1_3_AND2_NUM11 (.ZN (N573), .A1 (XNOR_1_1_AND2_NUM11_OUT), .A2 (XNOR_1_2_AND2_NUM11_OUT));
      wire XNOR_1_1_AND2_NUM12_OUT, XNOR_1_2_AND2_NUM12_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM12 (.ZN (XNOR_1_1_AND2_NUM12_OUT), .A1 (N1), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM12 (.ZN (XNOR_1_2_AND2_NUM12_OUT), .A1 (GND), .A2 (N460));
      NOR2_X1 XNOR_1_3_AND2_NUM12 (.ZN (N576), .A1 (XNOR_1_1_AND2_NUM12_OUT), .A2 (XNOR_1_2_AND2_NUM12_OUT));
      wire XNOR_1_1_AND2_NUM13_OUT, XNOR_1_2_AND2_NUM13_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM13 (.ZN (XNOR_1_1_AND2_NUM13_OUT), .A1 (N1), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM13 (.ZN (XNOR_1_2_AND2_NUM13_OUT), .A1 (GND), .A2 (N477));
      NOR2_X1 XNOR_1_3_AND2_NUM13 (.ZN (N579), .A1 (XNOR_1_1_AND2_NUM13_OUT), .A2 (XNOR_1_2_AND2_NUM13_OUT));
      wire XNOR_1_1_AND2_NUM14_OUT, XNOR_1_2_AND2_NUM14_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM14 (.ZN (XNOR_1_1_AND2_NUM14_OUT), .A1 (N1), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM14 (.ZN (XNOR_1_2_AND2_NUM14_OUT), .A1 (GND), .A2 (N494));
      NOR2_X1 XNOR_1_3_AND2_NUM14 (.ZN (N582), .A1 (XNOR_1_1_AND2_NUM14_OUT), .A2 (XNOR_1_2_AND2_NUM14_OUT));
      wire XNOR_1_1_AND2_NUM15_OUT, XNOR_1_2_AND2_NUM15_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM15 (.ZN (XNOR_1_1_AND2_NUM15_OUT), .A1 (N1), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM15 (.ZN (XNOR_1_2_AND2_NUM15_OUT), .A1 (GND), .A2 (N511));
      NOR2_X1 XNOR_1_3_AND2_NUM15 (.ZN (N585), .A1 (XNOR_1_1_AND2_NUM15_OUT), .A2 (XNOR_1_2_AND2_NUM15_OUT));
      wire XNOR_1_1_AND2_NUM16_OUT, XNOR_1_2_AND2_NUM16_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM16 (.ZN (XNOR_1_1_AND2_NUM16_OUT), .A1 (N1), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM16 (.ZN (XNOR_1_2_AND2_NUM16_OUT), .A1 (GND), .A2 (N528));
      NOR2_X1 XNOR_1_3_AND2_NUM16 (.ZN (N588), .A1 (XNOR_1_1_AND2_NUM16_OUT), .A2 (XNOR_1_2_AND2_NUM16_OUT));
      wire XNOR_1_1_AND2_NUM17_OUT, XNOR_1_2_AND2_NUM17_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM17 (.ZN (XNOR_1_1_AND2_NUM17_OUT), .A1 (N18), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM17 (.ZN (XNOR_1_2_AND2_NUM17_OUT), .A1 (GND), .A2 (N273));
      NOR2_X1 XNOR_1_3_AND2_NUM17 (.ZN (N591), .A1 (XNOR_1_1_AND2_NUM17_OUT), .A2 (XNOR_1_2_AND2_NUM17_OUT));
      wire XNOR_1_1_AND2_NUM18_OUT, XNOR_1_2_AND2_NUM18_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM18 (.ZN (XNOR_1_1_AND2_NUM18_OUT), .A1 (N18), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM18 (.ZN (XNOR_1_2_AND2_NUM18_OUT), .A1 (GND), .A2 (N290));
      NOR2_X1 XNOR_1_3_AND2_NUM18 (.ZN (N594), .A1 (XNOR_1_1_AND2_NUM18_OUT), .A2 (XNOR_1_2_AND2_NUM18_OUT));
      wire XNOR_1_1_AND2_NUM19_OUT, XNOR_1_2_AND2_NUM19_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM19 (.ZN (XNOR_1_1_AND2_NUM19_OUT), .A1 (N18), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM19 (.ZN (XNOR_1_2_AND2_NUM19_OUT), .A1 (GND), .A2 (N307));
      NOR2_X1 XNOR_1_3_AND2_NUM19 (.ZN (N597), .A1 (XNOR_1_1_AND2_NUM19_OUT), .A2 (XNOR_1_2_AND2_NUM19_OUT));
      wire XNOR_1_1_AND2_NUM20_OUT, XNOR_1_2_AND2_NUM20_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM20 (.ZN (XNOR_1_1_AND2_NUM20_OUT), .A1 (N18), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM20 (.ZN (XNOR_1_2_AND2_NUM20_OUT), .A1 (GND), .A2 (N324));
      NOR2_X1 XNOR_1_3_AND2_NUM20 (.ZN (N600), .A1 (XNOR_1_1_AND2_NUM20_OUT), .A2 (XNOR_1_2_AND2_NUM20_OUT));
      wire XNOR_1_1_AND2_NUM21_OUT, XNOR_1_2_AND2_NUM21_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM21 (.ZN (XNOR_1_1_AND2_NUM21_OUT), .A1 (N18), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM21 (.ZN (XNOR_1_2_AND2_NUM21_OUT), .A1 (GND), .A2 (N341));
      NOR2_X1 XNOR_1_3_AND2_NUM21 (.ZN (N603), .A1 (XNOR_1_1_AND2_NUM21_OUT), .A2 (XNOR_1_2_AND2_NUM21_OUT));
      wire XNOR_1_1_AND2_NUM22_OUT, XNOR_1_2_AND2_NUM22_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM22 (.ZN (XNOR_1_1_AND2_NUM22_OUT), .A1 (N18), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM22 (.ZN (XNOR_1_2_AND2_NUM22_OUT), .A1 (GND), .A2 (N358));
      NOR2_X1 XNOR_1_3_AND2_NUM22 (.ZN (N606), .A1 (XNOR_1_1_AND2_NUM22_OUT), .A2 (XNOR_1_2_AND2_NUM22_OUT));
      wire XNOR_1_1_AND2_NUM23_OUT, XNOR_1_2_AND2_NUM23_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM23 (.ZN (XNOR_1_1_AND2_NUM23_OUT), .A1 (N18), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM23 (.ZN (XNOR_1_2_AND2_NUM23_OUT), .A1 (GND), .A2 (N375));
      NOR2_X1 XNOR_1_3_AND2_NUM23 (.ZN (N609), .A1 (XNOR_1_1_AND2_NUM23_OUT), .A2 (XNOR_1_2_AND2_NUM23_OUT));
      wire XNOR_1_1_AND2_NUM24_OUT, XNOR_1_2_AND2_NUM24_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM24 (.ZN (XNOR_1_1_AND2_NUM24_OUT), .A1 (N18), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM24 (.ZN (XNOR_1_2_AND2_NUM24_OUT), .A1 (GND), .A2 (N392));
      NOR2_X1 XNOR_1_3_AND2_NUM24 (.ZN (N612), .A1 (XNOR_1_1_AND2_NUM24_OUT), .A2 (XNOR_1_2_AND2_NUM24_OUT));
      wire XNOR_1_1_AND2_NUM25_OUT, XNOR_1_2_AND2_NUM25_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM25 (.ZN (XNOR_1_1_AND2_NUM25_OUT), .A1 (N18), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM25 (.ZN (XNOR_1_2_AND2_NUM25_OUT), .A1 (GND), .A2 (N409));
      NOR2_X1 XNOR_1_3_AND2_NUM25 (.ZN (N615), .A1 (XNOR_1_1_AND2_NUM25_OUT), .A2 (XNOR_1_2_AND2_NUM25_OUT));
      wire XNOR_1_1_AND2_NUM26_OUT, XNOR_1_2_AND2_NUM26_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM26 (.ZN (XNOR_1_1_AND2_NUM26_OUT), .A1 (N18), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM26 (.ZN (XNOR_1_2_AND2_NUM26_OUT), .A1 (GND), .A2 (N426));
      NOR2_X1 XNOR_1_3_AND2_NUM26 (.ZN (N618), .A1 (XNOR_1_1_AND2_NUM26_OUT), .A2 (XNOR_1_2_AND2_NUM26_OUT));
      wire XNOR_1_1_AND2_NUM27_OUT, XNOR_1_2_AND2_NUM27_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM27 (.ZN (XNOR_1_1_AND2_NUM27_OUT), .A1 (N18), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM27 (.ZN (XNOR_1_2_AND2_NUM27_OUT), .A1 (GND), .A2 (N443));
      NOR2_X1 XNOR_1_3_AND2_NUM27 (.ZN (N621), .A1 (XNOR_1_1_AND2_NUM27_OUT), .A2 (XNOR_1_2_AND2_NUM27_OUT));
      wire XNOR_1_1_AND2_NUM28_OUT, XNOR_1_2_AND2_NUM28_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM28 (.ZN (XNOR_1_1_AND2_NUM28_OUT), .A1 (N18), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM28 (.ZN (XNOR_1_2_AND2_NUM28_OUT), .A1 (GND), .A2 (N460));
      NOR2_X1 XNOR_1_3_AND2_NUM28 (.ZN (N624), .A1 (XNOR_1_1_AND2_NUM28_OUT), .A2 (XNOR_1_2_AND2_NUM28_OUT));
      wire XNOR_1_1_AND2_NUM29_OUT, XNOR_1_2_AND2_NUM29_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM29 (.ZN (XNOR_1_1_AND2_NUM29_OUT), .A1 (N18), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM29 (.ZN (XNOR_1_2_AND2_NUM29_OUT), .A1 (GND), .A2 (N477));
      NOR2_X1 XNOR_1_3_AND2_NUM29 (.ZN (N627), .A1 (XNOR_1_1_AND2_NUM29_OUT), .A2 (XNOR_1_2_AND2_NUM29_OUT));
      wire XNOR_1_1_AND2_NUM30_OUT, XNOR_1_2_AND2_NUM30_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM30 (.ZN (XNOR_1_1_AND2_NUM30_OUT), .A1 (N18), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM30 (.ZN (XNOR_1_2_AND2_NUM30_OUT), .A1 (GND), .A2 (N494));
      NOR2_X1 XNOR_1_3_AND2_NUM30 (.ZN (N630), .A1 (XNOR_1_1_AND2_NUM30_OUT), .A2 (XNOR_1_2_AND2_NUM30_OUT));
      wire XNOR_1_1_AND2_NUM31_OUT, XNOR_1_2_AND2_NUM31_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM31 (.ZN (XNOR_1_1_AND2_NUM31_OUT), .A1 (N18), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM31 (.ZN (XNOR_1_2_AND2_NUM31_OUT), .A1 (GND), .A2 (N511));
      NOR2_X1 XNOR_1_3_AND2_NUM31 (.ZN (N633), .A1 (XNOR_1_1_AND2_NUM31_OUT), .A2 (XNOR_1_2_AND2_NUM31_OUT));
      wire XNOR_1_1_AND2_NUM32_OUT, XNOR_1_2_AND2_NUM32_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM32 (.ZN (XNOR_1_1_AND2_NUM32_OUT), .A1 (N18), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM32 (.ZN (XNOR_1_2_AND2_NUM32_OUT), .A1 (GND), .A2 (N528));
      NOR2_X1 XNOR_1_3_AND2_NUM32 (.ZN (N636), .A1 (XNOR_1_1_AND2_NUM32_OUT), .A2 (XNOR_1_2_AND2_NUM32_OUT));
      wire XNOR_1_1_AND2_NUM33_OUT, XNOR_1_2_AND2_NUM33_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM33 (.ZN (XNOR_1_1_AND2_NUM33_OUT), .A1 (N35), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM33 (.ZN (XNOR_1_2_AND2_NUM33_OUT), .A1 (GND), .A2 (N273));
      NOR2_X1 XNOR_1_3_AND2_NUM33 (.ZN (N639), .A1 (XNOR_1_1_AND2_NUM33_OUT), .A2 (XNOR_1_2_AND2_NUM33_OUT));
      wire XNOR_1_1_AND2_NUM34_OUT, XNOR_1_2_AND2_NUM34_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM34 (.ZN (XNOR_1_1_AND2_NUM34_OUT), .A1 (N35), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM34 (.ZN (XNOR_1_2_AND2_NUM34_OUT), .A1 (GND), .A2 (N290));
      NOR2_X1 XNOR_1_3_AND2_NUM34 (.ZN (N642), .A1 (XNOR_1_1_AND2_NUM34_OUT), .A2 (XNOR_1_2_AND2_NUM34_OUT));
      wire XNOR_1_1_AND2_NUM35_OUT, XNOR_1_2_AND2_NUM35_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM35 (.ZN (XNOR_1_1_AND2_NUM35_OUT), .A1 (N35), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM35 (.ZN (XNOR_1_2_AND2_NUM35_OUT), .A1 (GND), .A2 (N307));
      NOR2_X1 XNOR_1_3_AND2_NUM35 (.ZN (N645), .A1 (XNOR_1_1_AND2_NUM35_OUT), .A2 (XNOR_1_2_AND2_NUM35_OUT));
      wire XNOR_1_1_AND2_NUM36_OUT, XNOR_1_2_AND2_NUM36_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM36 (.ZN (XNOR_1_1_AND2_NUM36_OUT), .A1 (N35), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM36 (.ZN (XNOR_1_2_AND2_NUM36_OUT), .A1 (GND), .A2 (N324));
      NOR2_X1 XNOR_1_3_AND2_NUM36 (.ZN (N648), .A1 (XNOR_1_1_AND2_NUM36_OUT), .A2 (XNOR_1_2_AND2_NUM36_OUT));
      wire XNOR_1_1_AND2_NUM37_OUT, XNOR_1_2_AND2_NUM37_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM37 (.ZN (XNOR_1_1_AND2_NUM37_OUT), .A1 (N35), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM37 (.ZN (XNOR_1_2_AND2_NUM37_OUT), .A1 (GND), .A2 (N341));
      NOR2_X1 XNOR_1_3_AND2_NUM37 (.ZN (N651), .A1 (XNOR_1_1_AND2_NUM37_OUT), .A2 (XNOR_1_2_AND2_NUM37_OUT));
      wire XNOR_1_1_AND2_NUM38_OUT, XNOR_1_2_AND2_NUM38_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM38 (.ZN (XNOR_1_1_AND2_NUM38_OUT), .A1 (N35), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM38 (.ZN (XNOR_1_2_AND2_NUM38_OUT), .A1 (GND), .A2 (N358));
      NOR2_X1 XNOR_1_3_AND2_NUM38 (.ZN (N654), .A1 (XNOR_1_1_AND2_NUM38_OUT), .A2 (XNOR_1_2_AND2_NUM38_OUT));
      wire XNOR_1_1_AND2_NUM39_OUT, XNOR_1_2_AND2_NUM39_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM39 (.ZN (XNOR_1_1_AND2_NUM39_OUT), .A1 (N35), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM39 (.ZN (XNOR_1_2_AND2_NUM39_OUT), .A1 (GND), .A2 (N375));
      NOR2_X1 XNOR_1_3_AND2_NUM39 (.ZN (N657), .A1 (XNOR_1_1_AND2_NUM39_OUT), .A2 (XNOR_1_2_AND2_NUM39_OUT));
      wire XNOR_1_1_AND2_NUM40_OUT, XNOR_1_2_AND2_NUM40_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM40 (.ZN (XNOR_1_1_AND2_NUM40_OUT), .A1 (N35), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM40 (.ZN (XNOR_1_2_AND2_NUM40_OUT), .A1 (GND), .A2 (N392));
      NOR2_X1 XNOR_1_3_AND2_NUM40 (.ZN (N660), .A1 (XNOR_1_1_AND2_NUM40_OUT), .A2 (XNOR_1_2_AND2_NUM40_OUT));
      wire XNOR_1_1_AND2_NUM41_OUT, XNOR_1_2_AND2_NUM41_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM41 (.ZN (XNOR_1_1_AND2_NUM41_OUT), .A1 (N35), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM41 (.ZN (XNOR_1_2_AND2_NUM41_OUT), .A1 (GND), .A2 (N409));
      NOR2_X1 XNOR_1_3_AND2_NUM41 (.ZN (N663), .A1 (XNOR_1_1_AND2_NUM41_OUT), .A2 (XNOR_1_2_AND2_NUM41_OUT));
      wire XNOR_1_1_AND2_NUM42_OUT, XNOR_1_2_AND2_NUM42_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM42 (.ZN (XNOR_1_1_AND2_NUM42_OUT), .A1 (N35), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM42 (.ZN (XNOR_1_2_AND2_NUM42_OUT), .A1 (GND), .A2 (N426));
      NOR2_X1 XNOR_1_3_AND2_NUM42 (.ZN (N666), .A1 (XNOR_1_1_AND2_NUM42_OUT), .A2 (XNOR_1_2_AND2_NUM42_OUT));
      wire XNOR_1_1_AND2_NUM43_OUT, XNOR_1_2_AND2_NUM43_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM43 (.ZN (XNOR_1_1_AND2_NUM43_OUT), .A1 (N35), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM43 (.ZN (XNOR_1_2_AND2_NUM43_OUT), .A1 (GND), .A2 (N443));
      NOR2_X1 XNOR_1_3_AND2_NUM43 (.ZN (N669), .A1 (XNOR_1_1_AND2_NUM43_OUT), .A2 (XNOR_1_2_AND2_NUM43_OUT));
      wire XNOR_1_1_AND2_NUM44_OUT, XNOR_1_2_AND2_NUM44_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM44 (.ZN (XNOR_1_1_AND2_NUM44_OUT), .A1 (N35), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM44 (.ZN (XNOR_1_2_AND2_NUM44_OUT), .A1 (GND), .A2 (N460));
      NOR2_X1 XNOR_1_3_AND2_NUM44 (.ZN (N672), .A1 (XNOR_1_1_AND2_NUM44_OUT), .A2 (XNOR_1_2_AND2_NUM44_OUT));
      wire XNOR_1_1_AND2_NUM45_OUT, XNOR_1_2_AND2_NUM45_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM45 (.ZN (XNOR_1_1_AND2_NUM45_OUT), .A1 (N35), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM45 (.ZN (XNOR_1_2_AND2_NUM45_OUT), .A1 (GND), .A2 (N477));
      NOR2_X1 XNOR_1_3_AND2_NUM45 (.ZN (N675), .A1 (XNOR_1_1_AND2_NUM45_OUT), .A2 (XNOR_1_2_AND2_NUM45_OUT));
      wire XNOR_1_1_AND2_NUM46_OUT, XNOR_1_2_AND2_NUM46_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM46 (.ZN (XNOR_1_1_AND2_NUM46_OUT), .A1 (N35), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM46 (.ZN (XNOR_1_2_AND2_NUM46_OUT), .A1 (GND), .A2 (N494));
      NOR2_X1 XNOR_1_3_AND2_NUM46 (.ZN (N678), .A1 (XNOR_1_1_AND2_NUM46_OUT), .A2 (XNOR_1_2_AND2_NUM46_OUT));
      wire XNOR_1_1_AND2_NUM47_OUT, XNOR_1_2_AND2_NUM47_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM47 (.ZN (XNOR_1_1_AND2_NUM47_OUT), .A1 (N35), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM47 (.ZN (XNOR_1_2_AND2_NUM47_OUT), .A1 (GND), .A2 (N511));
      NOR2_X1 XNOR_1_3_AND2_NUM47 (.ZN (N681), .A1 (XNOR_1_1_AND2_NUM47_OUT), .A2 (XNOR_1_2_AND2_NUM47_OUT));
      wire XNOR_1_1_AND2_NUM48_OUT, XNOR_1_2_AND2_NUM48_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM48 (.ZN (XNOR_1_1_AND2_NUM48_OUT), .A1 (N35), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM48 (.ZN (XNOR_1_2_AND2_NUM48_OUT), .A1 (GND), .A2 (N528));
      NOR2_X1 XNOR_1_3_AND2_NUM48 (.ZN (N684), .A1 (XNOR_1_1_AND2_NUM48_OUT), .A2 (XNOR_1_2_AND2_NUM48_OUT));
      wire XNOR_1_1_AND2_NUM49_OUT, XNOR_1_2_AND2_NUM49_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM49 (.ZN (XNOR_1_1_AND2_NUM49_OUT), .A1 (N52), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM49 (.ZN (XNOR_1_2_AND2_NUM49_OUT), .A1 (GND), .A2 (N273));
      NOR2_X1 XNOR_1_3_AND2_NUM49 (.ZN (N687), .A1 (XNOR_1_1_AND2_NUM49_OUT), .A2 (XNOR_1_2_AND2_NUM49_OUT));
      wire XNOR_1_1_AND2_NUM50_OUT, XNOR_1_2_AND2_NUM50_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM50 (.ZN (XNOR_1_1_AND2_NUM50_OUT), .A1 (N52), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM50 (.ZN (XNOR_1_2_AND2_NUM50_OUT), .A1 (GND), .A2 (N290));
      NOR2_X1 XNOR_1_3_AND2_NUM50 (.ZN (N690), .A1 (XNOR_1_1_AND2_NUM50_OUT), .A2 (XNOR_1_2_AND2_NUM50_OUT));
      wire XNOR_1_1_AND2_NUM51_OUT, XNOR_1_2_AND2_NUM51_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM51 (.ZN (XNOR_1_1_AND2_NUM51_OUT), .A1 (N52), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM51 (.ZN (XNOR_1_2_AND2_NUM51_OUT), .A1 (GND), .A2 (N307));
      NOR2_X1 XNOR_1_3_AND2_NUM51 (.ZN (N693), .A1 (XNOR_1_1_AND2_NUM51_OUT), .A2 (XNOR_1_2_AND2_NUM51_OUT));
      wire XNOR_1_1_AND2_NUM52_OUT, XNOR_1_2_AND2_NUM52_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM52 (.ZN (XNOR_1_1_AND2_NUM52_OUT), .A1 (N52), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM52 (.ZN (XNOR_1_2_AND2_NUM52_OUT), .A1 (GND), .A2 (N324));
      NOR2_X1 XNOR_1_3_AND2_NUM52 (.ZN (N696), .A1 (XNOR_1_1_AND2_NUM52_OUT), .A2 (XNOR_1_2_AND2_NUM52_OUT));
      wire XNOR_1_1_AND2_NUM53_OUT, XNOR_1_2_AND2_NUM53_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM53 (.ZN (XNOR_1_1_AND2_NUM53_OUT), .A1 (N52), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM53 (.ZN (XNOR_1_2_AND2_NUM53_OUT), .A1 (GND), .A2 (N341));
      NOR2_X1 XNOR_1_3_AND2_NUM53 (.ZN (N699), .A1 (XNOR_1_1_AND2_NUM53_OUT), .A2 (XNOR_1_2_AND2_NUM53_OUT));
      wire XNOR_1_1_AND2_NUM54_OUT, XNOR_1_2_AND2_NUM54_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM54 (.ZN (XNOR_1_1_AND2_NUM54_OUT), .A1 (N52), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM54 (.ZN (XNOR_1_2_AND2_NUM54_OUT), .A1 (GND), .A2 (N358));
      NOR2_X1 XNOR_1_3_AND2_NUM54 (.ZN (N702), .A1 (XNOR_1_1_AND2_NUM54_OUT), .A2 (XNOR_1_2_AND2_NUM54_OUT));
      wire XNOR_1_1_AND2_NUM55_OUT, XNOR_1_2_AND2_NUM55_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM55 (.ZN (XNOR_1_1_AND2_NUM55_OUT), .A1 (N52), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM55 (.ZN (XNOR_1_2_AND2_NUM55_OUT), .A1 (GND), .A2 (N375));
      NOR2_X1 XNOR_1_3_AND2_NUM55 (.ZN (N705), .A1 (XNOR_1_1_AND2_NUM55_OUT), .A2 (XNOR_1_2_AND2_NUM55_OUT));
      wire XNOR_1_1_AND2_NUM56_OUT, XNOR_1_2_AND2_NUM56_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM56 (.ZN (XNOR_1_1_AND2_NUM56_OUT), .A1 (N52), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM56 (.ZN (XNOR_1_2_AND2_NUM56_OUT), .A1 (GND), .A2 (N392));
      NOR2_X1 XNOR_1_3_AND2_NUM56 (.ZN (N708), .A1 (XNOR_1_1_AND2_NUM56_OUT), .A2 (XNOR_1_2_AND2_NUM56_OUT));
      wire XNOR_1_1_AND2_NUM57_OUT, XNOR_1_2_AND2_NUM57_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM57 (.ZN (XNOR_1_1_AND2_NUM57_OUT), .A1 (N52), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM57 (.ZN (XNOR_1_2_AND2_NUM57_OUT), .A1 (GND), .A2 (N409));
      NOR2_X1 XNOR_1_3_AND2_NUM57 (.ZN (N711), .A1 (XNOR_1_1_AND2_NUM57_OUT), .A2 (XNOR_1_2_AND2_NUM57_OUT));
      wire XNOR_1_1_AND2_NUM58_OUT, XNOR_1_2_AND2_NUM58_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM58 (.ZN (XNOR_1_1_AND2_NUM58_OUT), .A1 (N52), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM58 (.ZN (XNOR_1_2_AND2_NUM58_OUT), .A1 (GND), .A2 (N426));
      NOR2_X1 XNOR_1_3_AND2_NUM58 (.ZN (N714), .A1 (XNOR_1_1_AND2_NUM58_OUT), .A2 (XNOR_1_2_AND2_NUM58_OUT));
      wire XNOR_1_1_AND2_NUM59_OUT, XNOR_1_2_AND2_NUM59_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM59 (.ZN (XNOR_1_1_AND2_NUM59_OUT), .A1 (N52), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM59 (.ZN (XNOR_1_2_AND2_NUM59_OUT), .A1 (GND), .A2 (N443));
      NOR2_X1 XNOR_1_3_AND2_NUM59 (.ZN (N717), .A1 (XNOR_1_1_AND2_NUM59_OUT), .A2 (XNOR_1_2_AND2_NUM59_OUT));
      wire XNOR_1_1_AND2_NUM60_OUT, XNOR_1_2_AND2_NUM60_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM60 (.ZN (XNOR_1_1_AND2_NUM60_OUT), .A1 (N52), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM60 (.ZN (XNOR_1_2_AND2_NUM60_OUT), .A1 (GND), .A2 (N460));
      NOR2_X1 XNOR_1_3_AND2_NUM60 (.ZN (N720), .A1 (XNOR_1_1_AND2_NUM60_OUT), .A2 (XNOR_1_2_AND2_NUM60_OUT));
      wire XNOR_1_1_AND2_NUM61_OUT, XNOR_1_2_AND2_NUM61_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM61 (.ZN (XNOR_1_1_AND2_NUM61_OUT), .A1 (N52), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM61 (.ZN (XNOR_1_2_AND2_NUM61_OUT), .A1 (GND), .A2 (N477));
      NOR2_X1 XNOR_1_3_AND2_NUM61 (.ZN (N723), .A1 (XNOR_1_1_AND2_NUM61_OUT), .A2 (XNOR_1_2_AND2_NUM61_OUT));
      wire XNOR_1_1_AND2_NUM62_OUT, XNOR_1_2_AND2_NUM62_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM62 (.ZN (XNOR_1_1_AND2_NUM62_OUT), .A1 (N52), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM62 (.ZN (XNOR_1_2_AND2_NUM62_OUT), .A1 (GND), .A2 (N494));
      NOR2_X1 XNOR_1_3_AND2_NUM62 (.ZN (N726), .A1 (XNOR_1_1_AND2_NUM62_OUT), .A2 (XNOR_1_2_AND2_NUM62_OUT));
      wire XNOR_1_1_AND2_NUM63_OUT, XNOR_1_2_AND2_NUM63_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM63 (.ZN (XNOR_1_1_AND2_NUM63_OUT), .A1 (N52), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM63 (.ZN (XNOR_1_2_AND2_NUM63_OUT), .A1 (GND), .A2 (N511));
      NOR2_X1 XNOR_1_3_AND2_NUM63 (.ZN (N729), .A1 (XNOR_1_1_AND2_NUM63_OUT), .A2 (XNOR_1_2_AND2_NUM63_OUT));
      wire XNOR_1_1_AND2_NUM64_OUT, XNOR_1_2_AND2_NUM64_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM64 (.ZN (XNOR_1_1_AND2_NUM64_OUT), .A1 (N52), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM64 (.ZN (XNOR_1_2_AND2_NUM64_OUT), .A1 (GND), .A2 (N528));
      NOR2_X1 XNOR_1_3_AND2_NUM64 (.ZN (N732), .A1 (XNOR_1_1_AND2_NUM64_OUT), .A2 (XNOR_1_2_AND2_NUM64_OUT));
      wire XNOR_1_1_AND2_NUM65_OUT, XNOR_1_2_AND2_NUM65_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM65 (.ZN (XNOR_1_1_AND2_NUM65_OUT), .A1 (N69), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM65 (.ZN (XNOR_1_2_AND2_NUM65_OUT), .A1 (GND), .A2 (N273));
      NOR2_X1 XNOR_1_3_AND2_NUM65 (.ZN (N735), .A1 (XNOR_1_1_AND2_NUM65_OUT), .A2 (XNOR_1_2_AND2_NUM65_OUT));
      wire XNOR_1_1_AND2_NUM66_OUT, XNOR_1_2_AND2_NUM66_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM66 (.ZN (XNOR_1_1_AND2_NUM66_OUT), .A1 (N69), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM66 (.ZN (XNOR_1_2_AND2_NUM66_OUT), .A1 (GND), .A2 (N290));
      NOR2_X1 XNOR_1_3_AND2_NUM66 (.ZN (N738), .A1 (XNOR_1_1_AND2_NUM66_OUT), .A2 (XNOR_1_2_AND2_NUM66_OUT));
      wire XNOR_1_1_AND2_NUM67_OUT, XNOR_1_2_AND2_NUM67_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM67 (.ZN (XNOR_1_1_AND2_NUM67_OUT), .A1 (N69), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM67 (.ZN (XNOR_1_2_AND2_NUM67_OUT), .A1 (GND), .A2 (N307));
      NOR2_X1 XNOR_1_3_AND2_NUM67 (.ZN (N741), .A1 (XNOR_1_1_AND2_NUM67_OUT), .A2 (XNOR_1_2_AND2_NUM67_OUT));
      wire XNOR_1_1_AND2_NUM68_OUT, XNOR_1_2_AND2_NUM68_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM68 (.ZN (XNOR_1_1_AND2_NUM68_OUT), .A1 (N69), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM68 (.ZN (XNOR_1_2_AND2_NUM68_OUT), .A1 (GND), .A2 (N324));
      NOR2_X1 XNOR_1_3_AND2_NUM68 (.ZN (N744), .A1 (XNOR_1_1_AND2_NUM68_OUT), .A2 (XNOR_1_2_AND2_NUM68_OUT));
      wire XNOR_1_1_AND2_NUM69_OUT, XNOR_1_2_AND2_NUM69_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM69 (.ZN (XNOR_1_1_AND2_NUM69_OUT), .A1 (N69), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM69 (.ZN (XNOR_1_2_AND2_NUM69_OUT), .A1 (GND), .A2 (N341));
      NOR2_X1 XNOR_1_3_AND2_NUM69 (.ZN (N747), .A1 (XNOR_1_1_AND2_NUM69_OUT), .A2 (XNOR_1_2_AND2_NUM69_OUT));
      wire XNOR_1_1_AND2_NUM70_OUT, XNOR_1_2_AND2_NUM70_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM70 (.ZN (XNOR_1_1_AND2_NUM70_OUT), .A1 (N69), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM70 (.ZN (XNOR_1_2_AND2_NUM70_OUT), .A1 (GND), .A2 (N358));
      NOR2_X1 XNOR_1_3_AND2_NUM70 (.ZN (N750), .A1 (XNOR_1_1_AND2_NUM70_OUT), .A2 (XNOR_1_2_AND2_NUM70_OUT));
      wire XNOR_1_1_AND2_NUM71_OUT, XNOR_1_2_AND2_NUM71_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM71 (.ZN (XNOR_1_1_AND2_NUM71_OUT), .A1 (N69), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM71 (.ZN (XNOR_1_2_AND2_NUM71_OUT), .A1 (GND), .A2 (N375));
      NOR2_X1 XNOR_1_3_AND2_NUM71 (.ZN (N753), .A1 (XNOR_1_1_AND2_NUM71_OUT), .A2 (XNOR_1_2_AND2_NUM71_OUT));
      wire XNOR_1_1_AND2_NUM72_OUT, XNOR_1_2_AND2_NUM72_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM72 (.ZN (XNOR_1_1_AND2_NUM72_OUT), .A1 (N69), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM72 (.ZN (XNOR_1_2_AND2_NUM72_OUT), .A1 (GND), .A2 (N392));
      NOR2_X1 XNOR_1_3_AND2_NUM72 (.ZN (N756), .A1 (XNOR_1_1_AND2_NUM72_OUT), .A2 (XNOR_1_2_AND2_NUM72_OUT));
      wire XNOR_1_1_AND2_NUM73_OUT, XNOR_1_2_AND2_NUM73_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM73 (.ZN (XNOR_1_1_AND2_NUM73_OUT), .A1 (N69), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM73 (.ZN (XNOR_1_2_AND2_NUM73_OUT), .A1 (GND), .A2 (N409));
      NOR2_X1 XNOR_1_3_AND2_NUM73 (.ZN (N759), .A1 (XNOR_1_1_AND2_NUM73_OUT), .A2 (XNOR_1_2_AND2_NUM73_OUT));
      wire XNOR_1_1_AND2_NUM74_OUT, XNOR_1_2_AND2_NUM74_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM74 (.ZN (XNOR_1_1_AND2_NUM74_OUT), .A1 (N69), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM74 (.ZN (XNOR_1_2_AND2_NUM74_OUT), .A1 (GND), .A2 (N426));
      NOR2_X1 XNOR_1_3_AND2_NUM74 (.ZN (N762), .A1 (XNOR_1_1_AND2_NUM74_OUT), .A2 (XNOR_1_2_AND2_NUM74_OUT));
      wire XNOR_1_1_AND2_NUM75_OUT, XNOR_1_2_AND2_NUM75_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM75 (.ZN (XNOR_1_1_AND2_NUM75_OUT), .A1 (N69), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM75 (.ZN (XNOR_1_2_AND2_NUM75_OUT), .A1 (GND), .A2 (N443));
      NOR2_X1 XNOR_1_3_AND2_NUM75 (.ZN (N765), .A1 (XNOR_1_1_AND2_NUM75_OUT), .A2 (XNOR_1_2_AND2_NUM75_OUT));
      wire XNOR_1_1_AND2_NUM76_OUT, XNOR_1_2_AND2_NUM76_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM76 (.ZN (XNOR_1_1_AND2_NUM76_OUT), .A1 (N69), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM76 (.ZN (XNOR_1_2_AND2_NUM76_OUT), .A1 (GND), .A2 (N460));
      NOR2_X1 XNOR_1_3_AND2_NUM76 (.ZN (N768), .A1 (XNOR_1_1_AND2_NUM76_OUT), .A2 (XNOR_1_2_AND2_NUM76_OUT));
      wire XNOR_1_1_AND2_NUM77_OUT, XNOR_1_2_AND2_NUM77_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM77 (.ZN (XNOR_1_1_AND2_NUM77_OUT), .A1 (N69), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM77 (.ZN (XNOR_1_2_AND2_NUM77_OUT), .A1 (GND), .A2 (N477));
      NOR2_X1 XNOR_1_3_AND2_NUM77 (.ZN (N771), .A1 (XNOR_1_1_AND2_NUM77_OUT), .A2 (XNOR_1_2_AND2_NUM77_OUT));
      wire XNOR_1_1_AND2_NUM78_OUT, XNOR_1_2_AND2_NUM78_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM78 (.ZN (XNOR_1_1_AND2_NUM78_OUT), .A1 (N69), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM78 (.ZN (XNOR_1_2_AND2_NUM78_OUT), .A1 (GND), .A2 (N494));
      NOR2_X1 XNOR_1_3_AND2_NUM78 (.ZN (N774), .A1 (XNOR_1_1_AND2_NUM78_OUT), .A2 (XNOR_1_2_AND2_NUM78_OUT));
      wire XNOR_1_1_AND2_NUM79_OUT, XNOR_1_2_AND2_NUM79_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM79 (.ZN (XNOR_1_1_AND2_NUM79_OUT), .A1 (N69), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM79 (.ZN (XNOR_1_2_AND2_NUM79_OUT), .A1 (GND), .A2 (N511));
      NOR2_X1 XNOR_1_3_AND2_NUM79 (.ZN (N777), .A1 (XNOR_1_1_AND2_NUM79_OUT), .A2 (XNOR_1_2_AND2_NUM79_OUT));
      wire XNOR_1_1_AND2_NUM80_OUT, XNOR_1_2_AND2_NUM80_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM80 (.ZN (XNOR_1_1_AND2_NUM80_OUT), .A1 (N69), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM80 (.ZN (XNOR_1_2_AND2_NUM80_OUT), .A1 (GND), .A2 (N528));
      NOR2_X1 XNOR_1_3_AND2_NUM80 (.ZN (N780), .A1 (XNOR_1_1_AND2_NUM80_OUT), .A2 (XNOR_1_2_AND2_NUM80_OUT));
      wire XNOR_1_1_AND2_NUM81_OUT, XNOR_1_2_AND2_NUM81_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM81 (.ZN (XNOR_1_1_AND2_NUM81_OUT), .A1 (N86), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM81 (.ZN (XNOR_1_2_AND2_NUM81_OUT), .A1 (GND), .A2 (N273));
      NOR2_X1 XNOR_1_3_AND2_NUM81 (.ZN (N783), .A1 (XNOR_1_1_AND2_NUM81_OUT), .A2 (XNOR_1_2_AND2_NUM81_OUT));
      wire XNOR_1_1_AND2_NUM82_OUT, XNOR_1_2_AND2_NUM82_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM82 (.ZN (XNOR_1_1_AND2_NUM82_OUT), .A1 (N86), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM82 (.ZN (XNOR_1_2_AND2_NUM82_OUT), .A1 (GND), .A2 (N290));
      NOR2_X1 XNOR_1_3_AND2_NUM82 (.ZN (N786), .A1 (XNOR_1_1_AND2_NUM82_OUT), .A2 (XNOR_1_2_AND2_NUM82_OUT));
      wire XNOR_1_1_AND2_NUM83_OUT, XNOR_1_2_AND2_NUM83_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM83 (.ZN (XNOR_1_1_AND2_NUM83_OUT), .A1 (N86), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM83 (.ZN (XNOR_1_2_AND2_NUM83_OUT), .A1 (GND), .A2 (N307));
      NOR2_X1 XNOR_1_3_AND2_NUM83 (.ZN (N789), .A1 (XNOR_1_1_AND2_NUM83_OUT), .A2 (XNOR_1_2_AND2_NUM83_OUT));
      wire XNOR_1_1_AND2_NUM84_OUT, XNOR_1_2_AND2_NUM84_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM84 (.ZN (XNOR_1_1_AND2_NUM84_OUT), .A1 (N86), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM84 (.ZN (XNOR_1_2_AND2_NUM84_OUT), .A1 (GND), .A2 (N324));
      NOR2_X1 XNOR_1_3_AND2_NUM84 (.ZN (N792), .A1 (XNOR_1_1_AND2_NUM84_OUT), .A2 (XNOR_1_2_AND2_NUM84_OUT));
      wire XNOR_1_1_AND2_NUM85_OUT, XNOR_1_2_AND2_NUM85_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM85 (.ZN (XNOR_1_1_AND2_NUM85_OUT), .A1 (N86), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM85 (.ZN (XNOR_1_2_AND2_NUM85_OUT), .A1 (GND), .A2 (N341));
      NOR2_X1 XNOR_1_3_AND2_NUM85 (.ZN (N795), .A1 (XNOR_1_1_AND2_NUM85_OUT), .A2 (XNOR_1_2_AND2_NUM85_OUT));
      wire XNOR_1_1_AND2_NUM86_OUT, XNOR_1_2_AND2_NUM86_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM86 (.ZN (XNOR_1_1_AND2_NUM86_OUT), .A1 (N86), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM86 (.ZN (XNOR_1_2_AND2_NUM86_OUT), .A1 (GND), .A2 (N358));
      NOR2_X1 XNOR_1_3_AND2_NUM86 (.ZN (N798), .A1 (XNOR_1_1_AND2_NUM86_OUT), .A2 (XNOR_1_2_AND2_NUM86_OUT));
      wire XNOR_1_1_AND2_NUM87_OUT, XNOR_1_2_AND2_NUM87_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM87 (.ZN (XNOR_1_1_AND2_NUM87_OUT), .A1 (N86), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM87 (.ZN (XNOR_1_2_AND2_NUM87_OUT), .A1 (GND), .A2 (N375));
      NOR2_X1 XNOR_1_3_AND2_NUM87 (.ZN (N801), .A1 (XNOR_1_1_AND2_NUM87_OUT), .A2 (XNOR_1_2_AND2_NUM87_OUT));
      wire XNOR_1_1_AND2_NUM88_OUT, XNOR_1_2_AND2_NUM88_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM88 (.ZN (XNOR_1_1_AND2_NUM88_OUT), .A1 (N86), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM88 (.ZN (XNOR_1_2_AND2_NUM88_OUT), .A1 (GND), .A2 (N392));
      NOR2_X1 XNOR_1_3_AND2_NUM88 (.ZN (N804), .A1 (XNOR_1_1_AND2_NUM88_OUT), .A2 (XNOR_1_2_AND2_NUM88_OUT));
      wire XNOR_1_1_AND2_NUM89_OUT, XNOR_1_2_AND2_NUM89_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM89 (.ZN (XNOR_1_1_AND2_NUM89_OUT), .A1 (N86), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM89 (.ZN (XNOR_1_2_AND2_NUM89_OUT), .A1 (GND), .A2 (N409));
      NOR2_X1 XNOR_1_3_AND2_NUM89 (.ZN (N807), .A1 (XNOR_1_1_AND2_NUM89_OUT), .A2 (XNOR_1_2_AND2_NUM89_OUT));
      wire XNOR_1_1_AND2_NUM90_OUT, XNOR_1_2_AND2_NUM90_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM90 (.ZN (XNOR_1_1_AND2_NUM90_OUT), .A1 (N86), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM90 (.ZN (XNOR_1_2_AND2_NUM90_OUT), .A1 (GND), .A2 (N426));
      NOR2_X1 XNOR_1_3_AND2_NUM90 (.ZN (N810), .A1 (XNOR_1_1_AND2_NUM90_OUT), .A2 (XNOR_1_2_AND2_NUM90_OUT));
      wire XNOR_1_1_AND2_NUM91_OUT, XNOR_1_2_AND2_NUM91_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM91 (.ZN (XNOR_1_1_AND2_NUM91_OUT), .A1 (N86), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM91 (.ZN (XNOR_1_2_AND2_NUM91_OUT), .A1 (GND), .A2 (N443));
      NOR2_X1 XNOR_1_3_AND2_NUM91 (.ZN (N813), .A1 (XNOR_1_1_AND2_NUM91_OUT), .A2 (XNOR_1_2_AND2_NUM91_OUT));
      wire XNOR_1_1_AND2_NUM92_OUT, XNOR_1_2_AND2_NUM92_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM92 (.ZN (XNOR_1_1_AND2_NUM92_OUT), .A1 (N86), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM92 (.ZN (XNOR_1_2_AND2_NUM92_OUT), .A1 (GND), .A2 (N460));
      NOR2_X1 XNOR_1_3_AND2_NUM92 (.ZN (N816), .A1 (XNOR_1_1_AND2_NUM92_OUT), .A2 (XNOR_1_2_AND2_NUM92_OUT));
      wire XNOR_1_1_AND2_NUM93_OUT, XNOR_1_2_AND2_NUM93_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM93 (.ZN (XNOR_1_1_AND2_NUM93_OUT), .A1 (N86), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM93 (.ZN (XNOR_1_2_AND2_NUM93_OUT), .A1 (GND), .A2 (N477));
      NOR2_X1 XNOR_1_3_AND2_NUM93 (.ZN (N819), .A1 (XNOR_1_1_AND2_NUM93_OUT), .A2 (XNOR_1_2_AND2_NUM93_OUT));
      wire XNOR_1_1_AND2_NUM94_OUT, XNOR_1_2_AND2_NUM94_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM94 (.ZN (XNOR_1_1_AND2_NUM94_OUT), .A1 (N86), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM94 (.ZN (XNOR_1_2_AND2_NUM94_OUT), .A1 (GND), .A2 (N494));
      NOR2_X1 XNOR_1_3_AND2_NUM94 (.ZN (N822), .A1 (XNOR_1_1_AND2_NUM94_OUT), .A2 (XNOR_1_2_AND2_NUM94_OUT));
      wire XNOR_1_1_AND2_NUM95_OUT, XNOR_1_2_AND2_NUM95_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM95 (.ZN (XNOR_1_1_AND2_NUM95_OUT), .A1 (N86), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM95 (.ZN (XNOR_1_2_AND2_NUM95_OUT), .A1 (GND), .A2 (N511));
      NOR2_X1 XNOR_1_3_AND2_NUM95 (.ZN (N825), .A1 (XNOR_1_1_AND2_NUM95_OUT), .A2 (XNOR_1_2_AND2_NUM95_OUT));
      wire XNOR_1_1_AND2_NUM96_OUT, XNOR_1_2_AND2_NUM96_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM96 (.ZN (XNOR_1_1_AND2_NUM96_OUT), .A1 (N86), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM96 (.ZN (XNOR_1_2_AND2_NUM96_OUT), .A1 (GND), .A2 (N528));
      NOR2_X1 XNOR_1_3_AND2_NUM96 (.ZN (N828), .A1 (XNOR_1_1_AND2_NUM96_OUT), .A2 (XNOR_1_2_AND2_NUM96_OUT));
      wire XNOR_1_1_AND2_NUM97_OUT, XNOR_1_2_AND2_NUM97_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM97 (.ZN (XNOR_1_1_AND2_NUM97_OUT), .A1 (N103), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM97 (.ZN (XNOR_1_2_AND2_NUM97_OUT), .A1 (GND), .A2 (N273));
      NOR2_X1 XNOR_1_3_AND2_NUM97 (.ZN (N831), .A1 (XNOR_1_1_AND2_NUM97_OUT), .A2 (XNOR_1_2_AND2_NUM97_OUT));
      wire XNOR_1_1_AND2_NUM98_OUT, XNOR_1_2_AND2_NUM98_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM98 (.ZN (XNOR_1_1_AND2_NUM98_OUT), .A1 (N103), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM98 (.ZN (XNOR_1_2_AND2_NUM98_OUT), .A1 (GND), .A2 (N290));
      NOR2_X1 XNOR_1_3_AND2_NUM98 (.ZN (N834), .A1 (XNOR_1_1_AND2_NUM98_OUT), .A2 (XNOR_1_2_AND2_NUM98_OUT));
      wire XNOR_1_1_AND2_NUM99_OUT, XNOR_1_2_AND2_NUM99_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM99 (.ZN (XNOR_1_1_AND2_NUM99_OUT), .A1 (N103), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM99 (.ZN (XNOR_1_2_AND2_NUM99_OUT), .A1 (GND), .A2 (N307));
      NOR2_X1 XNOR_1_3_AND2_NUM99 (.ZN (N837), .A1 (XNOR_1_1_AND2_NUM99_OUT), .A2 (XNOR_1_2_AND2_NUM99_OUT));
      wire XNOR_1_1_AND2_NUM100_OUT, XNOR_1_2_AND2_NUM100_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM100 (.ZN (XNOR_1_1_AND2_NUM100_OUT), .A1 (N103), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM100 (.ZN (XNOR_1_2_AND2_NUM100_OUT), .A1 (GND), .A2 (N324));
      NOR2_X1 XNOR_1_3_AND2_NUM100 (.ZN (N840), .A1 (XNOR_1_1_AND2_NUM100_OUT), .A2 (XNOR_1_2_AND2_NUM100_OUT));
      wire XNOR_1_1_AND2_NUM101_OUT, XNOR_1_2_AND2_NUM101_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM101 (.ZN (XNOR_1_1_AND2_NUM101_OUT), .A1 (N103), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM101 (.ZN (XNOR_1_2_AND2_NUM101_OUT), .A1 (GND), .A2 (N341));
      NOR2_X1 XNOR_1_3_AND2_NUM101 (.ZN (N843), .A1 (XNOR_1_1_AND2_NUM101_OUT), .A2 (XNOR_1_2_AND2_NUM101_OUT));
      wire XNOR_1_1_AND2_NUM102_OUT, XNOR_1_2_AND2_NUM102_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM102 (.ZN (XNOR_1_1_AND2_NUM102_OUT), .A1 (N103), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM102 (.ZN (XNOR_1_2_AND2_NUM102_OUT), .A1 (GND), .A2 (N358));
      NOR2_X1 XNOR_1_3_AND2_NUM102 (.ZN (N846), .A1 (XNOR_1_1_AND2_NUM102_OUT), .A2 (XNOR_1_2_AND2_NUM102_OUT));
      wire XNOR_1_1_AND2_NUM103_OUT, XNOR_1_2_AND2_NUM103_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM103 (.ZN (XNOR_1_1_AND2_NUM103_OUT), .A1 (N103), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM103 (.ZN (XNOR_1_2_AND2_NUM103_OUT), .A1 (GND), .A2 (N375));
      NOR2_X1 XNOR_1_3_AND2_NUM103 (.ZN (N849), .A1 (XNOR_1_1_AND2_NUM103_OUT), .A2 (XNOR_1_2_AND2_NUM103_OUT));
      wire XNOR_1_1_AND2_NUM104_OUT, XNOR_1_2_AND2_NUM104_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM104 (.ZN (XNOR_1_1_AND2_NUM104_OUT), .A1 (N103), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM104 (.ZN (XNOR_1_2_AND2_NUM104_OUT), .A1 (GND), .A2 (N392));
      NOR2_X1 XNOR_1_3_AND2_NUM104 (.ZN (N852), .A1 (XNOR_1_1_AND2_NUM104_OUT), .A2 (XNOR_1_2_AND2_NUM104_OUT));
      wire XNOR_1_1_AND2_NUM105_OUT, XNOR_1_2_AND2_NUM105_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM105 (.ZN (XNOR_1_1_AND2_NUM105_OUT), .A1 (N103), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM105 (.ZN (XNOR_1_2_AND2_NUM105_OUT), .A1 (GND), .A2 (N409));
      NOR2_X1 XNOR_1_3_AND2_NUM105 (.ZN (N855), .A1 (XNOR_1_1_AND2_NUM105_OUT), .A2 (XNOR_1_2_AND2_NUM105_OUT));
      wire XNOR_1_1_AND2_NUM106_OUT, XNOR_1_2_AND2_NUM106_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM106 (.ZN (XNOR_1_1_AND2_NUM106_OUT), .A1 (N103), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM106 (.ZN (XNOR_1_2_AND2_NUM106_OUT), .A1 (GND), .A2 (N426));
      NOR2_X1 XNOR_1_3_AND2_NUM106 (.ZN (N858), .A1 (XNOR_1_1_AND2_NUM106_OUT), .A2 (XNOR_1_2_AND2_NUM106_OUT));
      wire XNOR_1_1_AND2_NUM107_OUT, XNOR_1_2_AND2_NUM107_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM107 (.ZN (XNOR_1_1_AND2_NUM107_OUT), .A1 (N103), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM107 (.ZN (XNOR_1_2_AND2_NUM107_OUT), .A1 (GND), .A2 (N443));
      NOR2_X1 XNOR_1_3_AND2_NUM107 (.ZN (N861), .A1 (XNOR_1_1_AND2_NUM107_OUT), .A2 (XNOR_1_2_AND2_NUM107_OUT));
      wire XNOR_1_1_AND2_NUM108_OUT, XNOR_1_2_AND2_NUM108_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM108 (.ZN (XNOR_1_1_AND2_NUM108_OUT), .A1 (N103), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM108 (.ZN (XNOR_1_2_AND2_NUM108_OUT), .A1 (GND), .A2 (N460));
      NOR2_X1 XNOR_1_3_AND2_NUM108 (.ZN (N864), .A1 (XNOR_1_1_AND2_NUM108_OUT), .A2 (XNOR_1_2_AND2_NUM108_OUT));
      wire XNOR_1_1_AND2_NUM109_OUT, XNOR_1_2_AND2_NUM109_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM109 (.ZN (XNOR_1_1_AND2_NUM109_OUT), .A1 (N103), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM109 (.ZN (XNOR_1_2_AND2_NUM109_OUT), .A1 (GND), .A2 (N477));
      NOR2_X1 XNOR_1_3_AND2_NUM109 (.ZN (N867), .A1 (XNOR_1_1_AND2_NUM109_OUT), .A2 (XNOR_1_2_AND2_NUM109_OUT));
      wire XNOR_1_1_AND2_NUM110_OUT, XNOR_1_2_AND2_NUM110_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM110 (.ZN (XNOR_1_1_AND2_NUM110_OUT), .A1 (N103), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM110 (.ZN (XNOR_1_2_AND2_NUM110_OUT), .A1 (GND), .A2 (N494));
      NOR2_X1 XNOR_1_3_AND2_NUM110 (.ZN (N870), .A1 (XNOR_1_1_AND2_NUM110_OUT), .A2 (XNOR_1_2_AND2_NUM110_OUT));
      wire XNOR_1_1_AND2_NUM111_OUT, XNOR_1_2_AND2_NUM111_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM111 (.ZN (XNOR_1_1_AND2_NUM111_OUT), .A1 (N103), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM111 (.ZN (XNOR_1_2_AND2_NUM111_OUT), .A1 (GND), .A2 (N511));
      NOR2_X1 XNOR_1_3_AND2_NUM111 (.ZN (N873), .A1 (XNOR_1_1_AND2_NUM111_OUT), .A2 (XNOR_1_2_AND2_NUM111_OUT));
      wire XNOR_1_1_AND2_NUM112_OUT, XNOR_1_2_AND2_NUM112_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM112 (.ZN (XNOR_1_1_AND2_NUM112_OUT), .A1 (N103), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM112 (.ZN (XNOR_1_2_AND2_NUM112_OUT), .A1 (GND), .A2 (N528));
      NOR2_X1 XNOR_1_3_AND2_NUM112 (.ZN (N876), .A1 (XNOR_1_1_AND2_NUM112_OUT), .A2 (XNOR_1_2_AND2_NUM112_OUT));
      wire XNOR_1_1_AND2_NUM113_OUT, XNOR_1_2_AND2_NUM113_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM113 (.ZN (XNOR_1_1_AND2_NUM113_OUT), .A1 (N120), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM113 (.ZN (XNOR_1_2_AND2_NUM113_OUT), .A1 (GND), .A2 (N273));
      NOR2_X1 XNOR_1_3_AND2_NUM113 (.ZN (N879), .A1 (XNOR_1_1_AND2_NUM113_OUT), .A2 (XNOR_1_2_AND2_NUM113_OUT));
      wire XNOR_1_1_AND2_NUM114_OUT, XNOR_1_2_AND2_NUM114_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM114 (.ZN (XNOR_1_1_AND2_NUM114_OUT), .A1 (N120), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM114 (.ZN (XNOR_1_2_AND2_NUM114_OUT), .A1 (GND), .A2 (N290));
      NOR2_X1 XNOR_1_3_AND2_NUM114 (.ZN (N882), .A1 (XNOR_1_1_AND2_NUM114_OUT), .A2 (XNOR_1_2_AND2_NUM114_OUT));
      wire XNOR_1_1_AND2_NUM115_OUT, XNOR_1_2_AND2_NUM115_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM115 (.ZN (XNOR_1_1_AND2_NUM115_OUT), .A1 (N120), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM115 (.ZN (XNOR_1_2_AND2_NUM115_OUT), .A1 (GND), .A2 (N307));
      NOR2_X1 XNOR_1_3_AND2_NUM115 (.ZN (N885), .A1 (XNOR_1_1_AND2_NUM115_OUT), .A2 (XNOR_1_2_AND2_NUM115_OUT));
      wire XNOR_1_1_AND2_NUM116_OUT, XNOR_1_2_AND2_NUM116_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM116 (.ZN (XNOR_1_1_AND2_NUM116_OUT), .A1 (N120), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM116 (.ZN (XNOR_1_2_AND2_NUM116_OUT), .A1 (GND), .A2 (N324));
      NOR2_X1 XNOR_1_3_AND2_NUM116 (.ZN (N888), .A1 (XNOR_1_1_AND2_NUM116_OUT), .A2 (XNOR_1_2_AND2_NUM116_OUT));
      wire XNOR_1_1_AND2_NUM117_OUT, XNOR_1_2_AND2_NUM117_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM117 (.ZN (XNOR_1_1_AND2_NUM117_OUT), .A1 (N120), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM117 (.ZN (XNOR_1_2_AND2_NUM117_OUT), .A1 (GND), .A2 (N341));
      NOR2_X1 XNOR_1_3_AND2_NUM117 (.ZN (N891), .A1 (XNOR_1_1_AND2_NUM117_OUT), .A2 (XNOR_1_2_AND2_NUM117_OUT));
      wire XNOR_1_1_AND2_NUM118_OUT, XNOR_1_2_AND2_NUM118_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM118 (.ZN (XNOR_1_1_AND2_NUM118_OUT), .A1 (N120), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM118 (.ZN (XNOR_1_2_AND2_NUM118_OUT), .A1 (GND), .A2 (N358));
      NOR2_X1 XNOR_1_3_AND2_NUM118 (.ZN (N894), .A1 (XNOR_1_1_AND2_NUM118_OUT), .A2 (XNOR_1_2_AND2_NUM118_OUT));
      wire XNOR_1_1_AND2_NUM119_OUT, XNOR_1_2_AND2_NUM119_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM119 (.ZN (XNOR_1_1_AND2_NUM119_OUT), .A1 (N120), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM119 (.ZN (XNOR_1_2_AND2_NUM119_OUT), .A1 (GND), .A2 (N375));
      NOR2_X1 XNOR_1_3_AND2_NUM119 (.ZN (N897), .A1 (XNOR_1_1_AND2_NUM119_OUT), .A2 (XNOR_1_2_AND2_NUM119_OUT));
      wire XNOR_1_1_AND2_NUM120_OUT, XNOR_1_2_AND2_NUM120_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM120 (.ZN (XNOR_1_1_AND2_NUM120_OUT), .A1 (N120), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM120 (.ZN (XNOR_1_2_AND2_NUM120_OUT), .A1 (GND), .A2 (N392));
      NOR2_X1 XNOR_1_3_AND2_NUM120 (.ZN (N900), .A1 (XNOR_1_1_AND2_NUM120_OUT), .A2 (XNOR_1_2_AND2_NUM120_OUT));
      wire XNOR_1_1_AND2_NUM121_OUT, XNOR_1_2_AND2_NUM121_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM121 (.ZN (XNOR_1_1_AND2_NUM121_OUT), .A1 (N120), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM121 (.ZN (XNOR_1_2_AND2_NUM121_OUT), .A1 (GND), .A2 (N409));
      NOR2_X1 XNOR_1_3_AND2_NUM121 (.ZN (N903), .A1 (XNOR_1_1_AND2_NUM121_OUT), .A2 (XNOR_1_2_AND2_NUM121_OUT));
      wire XNOR_1_1_AND2_NUM122_OUT, XNOR_1_2_AND2_NUM122_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM122 (.ZN (XNOR_1_1_AND2_NUM122_OUT), .A1 (N120), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM122 (.ZN (XNOR_1_2_AND2_NUM122_OUT), .A1 (GND), .A2 (N426));
      NOR2_X1 XNOR_1_3_AND2_NUM122 (.ZN (N906), .A1 (XNOR_1_1_AND2_NUM122_OUT), .A2 (XNOR_1_2_AND2_NUM122_OUT));
      wire XNOR_1_1_AND2_NUM123_OUT, XNOR_1_2_AND2_NUM123_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM123 (.ZN (XNOR_1_1_AND2_NUM123_OUT), .A1 (N120), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM123 (.ZN (XNOR_1_2_AND2_NUM123_OUT), .A1 (GND), .A2 (N443));
      NOR2_X1 XNOR_1_3_AND2_NUM123 (.ZN (N909), .A1 (XNOR_1_1_AND2_NUM123_OUT), .A2 (XNOR_1_2_AND2_NUM123_OUT));
      wire XNOR_1_1_AND2_NUM124_OUT, XNOR_1_2_AND2_NUM124_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM124 (.ZN (XNOR_1_1_AND2_NUM124_OUT), .A1 (N120), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM124 (.ZN (XNOR_1_2_AND2_NUM124_OUT), .A1 (GND), .A2 (N460));
      NOR2_X1 XNOR_1_3_AND2_NUM124 (.ZN (N912), .A1 (XNOR_1_1_AND2_NUM124_OUT), .A2 (XNOR_1_2_AND2_NUM124_OUT));
      wire XNOR_1_1_AND2_NUM125_OUT, XNOR_1_2_AND2_NUM125_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM125 (.ZN (XNOR_1_1_AND2_NUM125_OUT), .A1 (N120), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM125 (.ZN (XNOR_1_2_AND2_NUM125_OUT), .A1 (GND), .A2 (N477));
      NOR2_X1 XNOR_1_3_AND2_NUM125 (.ZN (N915), .A1 (XNOR_1_1_AND2_NUM125_OUT), .A2 (XNOR_1_2_AND2_NUM125_OUT));
      wire XNOR_1_1_AND2_NUM126_OUT, XNOR_1_2_AND2_NUM126_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM126 (.ZN (XNOR_1_1_AND2_NUM126_OUT), .A1 (N120), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM126 (.ZN (XNOR_1_2_AND2_NUM126_OUT), .A1 (GND), .A2 (N494));
      NOR2_X1 XNOR_1_3_AND2_NUM126 (.ZN (N918), .A1 (XNOR_1_1_AND2_NUM126_OUT), .A2 (XNOR_1_2_AND2_NUM126_OUT));
      wire XNOR_1_1_AND2_NUM127_OUT, XNOR_1_2_AND2_NUM127_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM127 (.ZN (XNOR_1_1_AND2_NUM127_OUT), .A1 (N120), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM127 (.ZN (XNOR_1_2_AND2_NUM127_OUT), .A1 (GND), .A2 (N511));
      NOR2_X1 XNOR_1_3_AND2_NUM127 (.ZN (N921), .A1 (XNOR_1_1_AND2_NUM127_OUT), .A2 (XNOR_1_2_AND2_NUM127_OUT));
      wire XNOR_1_1_AND2_NUM128_OUT, XNOR_1_2_AND2_NUM128_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM128 (.ZN (XNOR_1_1_AND2_NUM128_OUT), .A1 (N120), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM128 (.ZN (XNOR_1_2_AND2_NUM128_OUT), .A1 (GND), .A2 (N528));
      NOR2_X1 XNOR_1_3_AND2_NUM128 (.ZN (N924), .A1 (XNOR_1_1_AND2_NUM128_OUT), .A2 (XNOR_1_2_AND2_NUM128_OUT));
      wire XNOR_1_1_AND2_NUM129_OUT, XNOR_1_2_AND2_NUM129_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM129 (.ZN (XNOR_1_1_AND2_NUM129_OUT), .A1 (N137), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM129 (.ZN (XNOR_1_2_AND2_NUM129_OUT), .A1 (GND), .A2 (N273));
      NOR2_X1 XNOR_1_3_AND2_NUM129 (.ZN (N927), .A1 (XNOR_1_1_AND2_NUM129_OUT), .A2 (XNOR_1_2_AND2_NUM129_OUT));
      wire XNOR_1_1_AND2_NUM130_OUT, XNOR_1_2_AND2_NUM130_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM130 (.ZN (XNOR_1_1_AND2_NUM130_OUT), .A1 (N137), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM130 (.ZN (XNOR_1_2_AND2_NUM130_OUT), .A1 (GND), .A2 (N290));
      NOR2_X1 XNOR_1_3_AND2_NUM130 (.ZN (N930), .A1 (XNOR_1_1_AND2_NUM130_OUT), .A2 (XNOR_1_2_AND2_NUM130_OUT));
      wire XNOR_1_1_AND2_NUM131_OUT, XNOR_1_2_AND2_NUM131_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM131 (.ZN (XNOR_1_1_AND2_NUM131_OUT), .A1 (N137), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM131 (.ZN (XNOR_1_2_AND2_NUM131_OUT), .A1 (GND), .A2 (N307));
      NOR2_X1 XNOR_1_3_AND2_NUM131 (.ZN (N933), .A1 (XNOR_1_1_AND2_NUM131_OUT), .A2 (XNOR_1_2_AND2_NUM131_OUT));
      wire XNOR_1_1_AND2_NUM132_OUT, XNOR_1_2_AND2_NUM132_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM132 (.ZN (XNOR_1_1_AND2_NUM132_OUT), .A1 (N137), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM132 (.ZN (XNOR_1_2_AND2_NUM132_OUT), .A1 (GND), .A2 (N324));
      NOR2_X1 XNOR_1_3_AND2_NUM132 (.ZN (N936), .A1 (XNOR_1_1_AND2_NUM132_OUT), .A2 (XNOR_1_2_AND2_NUM132_OUT));
      wire XNOR_1_1_AND2_NUM133_OUT, XNOR_1_2_AND2_NUM133_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM133 (.ZN (XNOR_1_1_AND2_NUM133_OUT), .A1 (N137), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM133 (.ZN (XNOR_1_2_AND2_NUM133_OUT), .A1 (GND), .A2 (N341));
      NOR2_X1 XNOR_1_3_AND2_NUM133 (.ZN (N939), .A1 (XNOR_1_1_AND2_NUM133_OUT), .A2 (XNOR_1_2_AND2_NUM133_OUT));
      wire XNOR_1_1_AND2_NUM134_OUT, XNOR_1_2_AND2_NUM134_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM134 (.ZN (XNOR_1_1_AND2_NUM134_OUT), .A1 (N137), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM134 (.ZN (XNOR_1_2_AND2_NUM134_OUT), .A1 (GND), .A2 (N358));
      NOR2_X1 XNOR_1_3_AND2_NUM134 (.ZN (N942), .A1 (XNOR_1_1_AND2_NUM134_OUT), .A2 (XNOR_1_2_AND2_NUM134_OUT));
      wire XNOR_1_1_AND2_NUM135_OUT, XNOR_1_2_AND2_NUM135_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM135 (.ZN (XNOR_1_1_AND2_NUM135_OUT), .A1 (N137), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM135 (.ZN (XNOR_1_2_AND2_NUM135_OUT), .A1 (GND), .A2 (N375));
      NOR2_X1 XNOR_1_3_AND2_NUM135 (.ZN (N945), .A1 (XNOR_1_1_AND2_NUM135_OUT), .A2 (XNOR_1_2_AND2_NUM135_OUT));
      wire XNOR_1_1_AND2_NUM136_OUT, XNOR_1_2_AND2_NUM136_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM136 (.ZN (XNOR_1_1_AND2_NUM136_OUT), .A1 (N137), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM136 (.ZN (XNOR_1_2_AND2_NUM136_OUT), .A1 (GND), .A2 (N392));
      NOR2_X1 XNOR_1_3_AND2_NUM136 (.ZN (N948), .A1 (XNOR_1_1_AND2_NUM136_OUT), .A2 (XNOR_1_2_AND2_NUM136_OUT));
      wire XNOR_1_1_AND2_NUM137_OUT, XNOR_1_2_AND2_NUM137_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM137 (.ZN (XNOR_1_1_AND2_NUM137_OUT), .A1 (N137), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM137 (.ZN (XNOR_1_2_AND2_NUM137_OUT), .A1 (GND), .A2 (N409));
      NOR2_X1 XNOR_1_3_AND2_NUM137 (.ZN (N951), .A1 (XNOR_1_1_AND2_NUM137_OUT), .A2 (XNOR_1_2_AND2_NUM137_OUT));
      wire XNOR_1_1_AND2_NUM138_OUT, XNOR_1_2_AND2_NUM138_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM138 (.ZN (XNOR_1_1_AND2_NUM138_OUT), .A1 (N137), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM138 (.ZN (XNOR_1_2_AND2_NUM138_OUT), .A1 (GND), .A2 (N426));
      NOR2_X1 XNOR_1_3_AND2_NUM138 (.ZN (N954), .A1 (XNOR_1_1_AND2_NUM138_OUT), .A2 (XNOR_1_2_AND2_NUM138_OUT));
      wire XNOR_1_1_AND2_NUM139_OUT, XNOR_1_2_AND2_NUM139_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM139 (.ZN (XNOR_1_1_AND2_NUM139_OUT), .A1 (N137), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM139 (.ZN (XNOR_1_2_AND2_NUM139_OUT), .A1 (GND), .A2 (N443));
      NOR2_X1 XNOR_1_3_AND2_NUM139 (.ZN (N957), .A1 (XNOR_1_1_AND2_NUM139_OUT), .A2 (XNOR_1_2_AND2_NUM139_OUT));
      wire XNOR_1_1_AND2_NUM140_OUT, XNOR_1_2_AND2_NUM140_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM140 (.ZN (XNOR_1_1_AND2_NUM140_OUT), .A1 (N137), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM140 (.ZN (XNOR_1_2_AND2_NUM140_OUT), .A1 (GND), .A2 (N460));
      NOR2_X1 XNOR_1_3_AND2_NUM140 (.ZN (N960), .A1 (XNOR_1_1_AND2_NUM140_OUT), .A2 (XNOR_1_2_AND2_NUM140_OUT));
      wire XNOR_1_1_AND2_NUM141_OUT, XNOR_1_2_AND2_NUM141_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM141 (.ZN (XNOR_1_1_AND2_NUM141_OUT), .A1 (N137), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM141 (.ZN (XNOR_1_2_AND2_NUM141_OUT), .A1 (GND), .A2 (N477));
      NOR2_X1 XNOR_1_3_AND2_NUM141 (.ZN (N963), .A1 (XNOR_1_1_AND2_NUM141_OUT), .A2 (XNOR_1_2_AND2_NUM141_OUT));
      wire XNOR_1_1_AND2_NUM142_OUT, XNOR_1_2_AND2_NUM142_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM142 (.ZN (XNOR_1_1_AND2_NUM142_OUT), .A1 (N137), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM142 (.ZN (XNOR_1_2_AND2_NUM142_OUT), .A1 (GND), .A2 (N494));
      NOR2_X1 XNOR_1_3_AND2_NUM142 (.ZN (N966), .A1 (XNOR_1_1_AND2_NUM142_OUT), .A2 (XNOR_1_2_AND2_NUM142_OUT));
      wire XNOR_1_1_AND2_NUM143_OUT, XNOR_1_2_AND2_NUM143_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM143 (.ZN (XNOR_1_1_AND2_NUM143_OUT), .A1 (N137), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM143 (.ZN (XNOR_1_2_AND2_NUM143_OUT), .A1 (GND), .A2 (N511));
      NOR2_X1 XNOR_1_3_AND2_NUM143 (.ZN (N969), .A1 (XNOR_1_1_AND2_NUM143_OUT), .A2 (XNOR_1_2_AND2_NUM143_OUT));
      wire XNOR_1_1_AND2_NUM144_OUT, XNOR_1_2_AND2_NUM144_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM144 (.ZN (XNOR_1_1_AND2_NUM144_OUT), .A1 (N137), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM144 (.ZN (XNOR_1_2_AND2_NUM144_OUT), .A1 (GND), .A2 (N528));
      NOR2_X1 XNOR_1_3_AND2_NUM144 (.ZN (N972), .A1 (XNOR_1_1_AND2_NUM144_OUT), .A2 (XNOR_1_2_AND2_NUM144_OUT));
      wire XNOR_1_1_AND2_NUM145_OUT, XNOR_1_2_AND2_NUM145_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM145 (.ZN (XNOR_1_1_AND2_NUM145_OUT), .A1 (N154), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM145 (.ZN (XNOR_1_2_AND2_NUM145_OUT), .A1 (GND), .A2 (N273));
      NOR2_X1 XNOR_1_3_AND2_NUM145 (.ZN (N975), .A1 (XNOR_1_1_AND2_NUM145_OUT), .A2 (XNOR_1_2_AND2_NUM145_OUT));
      wire XNOR_1_1_AND2_NUM146_OUT, XNOR_1_2_AND2_NUM146_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM146 (.ZN (XNOR_1_1_AND2_NUM146_OUT), .A1 (N154), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM146 (.ZN (XNOR_1_2_AND2_NUM146_OUT), .A1 (GND), .A2 (N290));
      NOR2_X1 XNOR_1_3_AND2_NUM146 (.ZN (N978), .A1 (XNOR_1_1_AND2_NUM146_OUT), .A2 (XNOR_1_2_AND2_NUM146_OUT));
      wire XNOR_1_1_AND2_NUM147_OUT, XNOR_1_2_AND2_NUM147_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM147 (.ZN (XNOR_1_1_AND2_NUM147_OUT), .A1 (N154), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM147 (.ZN (XNOR_1_2_AND2_NUM147_OUT), .A1 (GND), .A2 (N307));
      NOR2_X1 XNOR_1_3_AND2_NUM147 (.ZN (N981), .A1 (XNOR_1_1_AND2_NUM147_OUT), .A2 (XNOR_1_2_AND2_NUM147_OUT));
      wire XNOR_1_1_AND2_NUM148_OUT, XNOR_1_2_AND2_NUM148_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM148 (.ZN (XNOR_1_1_AND2_NUM148_OUT), .A1 (N154), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM148 (.ZN (XNOR_1_2_AND2_NUM148_OUT), .A1 (GND), .A2 (N324));
      NOR2_X1 XNOR_1_3_AND2_NUM148 (.ZN (N984), .A1 (XNOR_1_1_AND2_NUM148_OUT), .A2 (XNOR_1_2_AND2_NUM148_OUT));
      wire XNOR_1_1_AND2_NUM149_OUT, XNOR_1_2_AND2_NUM149_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM149 (.ZN (XNOR_1_1_AND2_NUM149_OUT), .A1 (N154), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM149 (.ZN (XNOR_1_2_AND2_NUM149_OUT), .A1 (GND), .A2 (N341));
      NOR2_X1 XNOR_1_3_AND2_NUM149 (.ZN (N987), .A1 (XNOR_1_1_AND2_NUM149_OUT), .A2 (XNOR_1_2_AND2_NUM149_OUT));
      wire XNOR_1_1_AND2_NUM150_OUT, XNOR_1_2_AND2_NUM150_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM150 (.ZN (XNOR_1_1_AND2_NUM150_OUT), .A1 (N154), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM150 (.ZN (XNOR_1_2_AND2_NUM150_OUT), .A1 (GND), .A2 (N358));
      NOR2_X1 XNOR_1_3_AND2_NUM150 (.ZN (N990), .A1 (XNOR_1_1_AND2_NUM150_OUT), .A2 (XNOR_1_2_AND2_NUM150_OUT));
      wire XNOR_1_1_AND2_NUM151_OUT, XNOR_1_2_AND2_NUM151_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM151 (.ZN (XNOR_1_1_AND2_NUM151_OUT), .A1 (N154), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM151 (.ZN (XNOR_1_2_AND2_NUM151_OUT), .A1 (GND), .A2 (N375));
      NOR2_X1 XNOR_1_3_AND2_NUM151 (.ZN (N993), .A1 (XNOR_1_1_AND2_NUM151_OUT), .A2 (XNOR_1_2_AND2_NUM151_OUT));
      wire XNOR_1_1_AND2_NUM152_OUT, XNOR_1_2_AND2_NUM152_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM152 (.ZN (XNOR_1_1_AND2_NUM152_OUT), .A1 (N154), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM152 (.ZN (XNOR_1_2_AND2_NUM152_OUT), .A1 (GND), .A2 (N392));
      NOR2_X1 XNOR_1_3_AND2_NUM152 (.ZN (N996), .A1 (XNOR_1_1_AND2_NUM152_OUT), .A2 (XNOR_1_2_AND2_NUM152_OUT));
      wire XNOR_1_1_AND2_NUM153_OUT, XNOR_1_2_AND2_NUM153_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM153 (.ZN (XNOR_1_1_AND2_NUM153_OUT), .A1 (N154), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM153 (.ZN (XNOR_1_2_AND2_NUM153_OUT), .A1 (GND), .A2 (N409));
      NOR2_X1 XNOR_1_3_AND2_NUM153 (.ZN (N999), .A1 (XNOR_1_1_AND2_NUM153_OUT), .A2 (XNOR_1_2_AND2_NUM153_OUT));
      wire XNOR_1_1_AND2_NUM154_OUT, XNOR_1_2_AND2_NUM154_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM154 (.ZN (XNOR_1_1_AND2_NUM154_OUT), .A1 (N154), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM154 (.ZN (XNOR_1_2_AND2_NUM154_OUT), .A1 (GND), .A2 (N426));
      NOR2_X1 XNOR_1_3_AND2_NUM154 (.ZN (N1002), .A1 (XNOR_1_1_AND2_NUM154_OUT), .A2 (XNOR_1_2_AND2_NUM154_OUT));
      wire XNOR_1_1_AND2_NUM155_OUT, XNOR_1_2_AND2_NUM155_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM155 (.ZN (XNOR_1_1_AND2_NUM155_OUT), .A1 (N154), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM155 (.ZN (XNOR_1_2_AND2_NUM155_OUT), .A1 (GND), .A2 (N443));
      NOR2_X1 XNOR_1_3_AND2_NUM155 (.ZN (N1005), .A1 (XNOR_1_1_AND2_NUM155_OUT), .A2 (XNOR_1_2_AND2_NUM155_OUT));
      wire XNOR_1_1_AND2_NUM156_OUT, XNOR_1_2_AND2_NUM156_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM156 (.ZN (XNOR_1_1_AND2_NUM156_OUT), .A1 (N154), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM156 (.ZN (XNOR_1_2_AND2_NUM156_OUT), .A1 (GND), .A2 (N460));
      NOR2_X1 XNOR_1_3_AND2_NUM156 (.ZN (N1008), .A1 (XNOR_1_1_AND2_NUM156_OUT), .A2 (XNOR_1_2_AND2_NUM156_OUT));
      wire XNOR_1_1_AND2_NUM157_OUT, XNOR_1_2_AND2_NUM157_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM157 (.ZN (XNOR_1_1_AND2_NUM157_OUT), .A1 (N154), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM157 (.ZN (XNOR_1_2_AND2_NUM157_OUT), .A1 (GND), .A2 (N477));
      NOR2_X1 XNOR_1_3_AND2_NUM157 (.ZN (N1011), .A1 (XNOR_1_1_AND2_NUM157_OUT), .A2 (XNOR_1_2_AND2_NUM157_OUT));
      wire XNOR_1_1_AND2_NUM158_OUT, XNOR_1_2_AND2_NUM158_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM158 (.ZN (XNOR_1_1_AND2_NUM158_OUT), .A1 (N154), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM158 (.ZN (XNOR_1_2_AND2_NUM158_OUT), .A1 (GND), .A2 (N494));
      NOR2_X1 XNOR_1_3_AND2_NUM158 (.ZN (N1014), .A1 (XNOR_1_1_AND2_NUM158_OUT), .A2 (XNOR_1_2_AND2_NUM158_OUT));
      wire XNOR_1_1_AND2_NUM159_OUT, XNOR_1_2_AND2_NUM159_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM159 (.ZN (XNOR_1_1_AND2_NUM159_OUT), .A1 (N154), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM159 (.ZN (XNOR_1_2_AND2_NUM159_OUT), .A1 (GND), .A2 (N511));
      NOR2_X1 XNOR_1_3_AND2_NUM159 (.ZN (N1017), .A1 (XNOR_1_1_AND2_NUM159_OUT), .A2 (XNOR_1_2_AND2_NUM159_OUT));
      wire XNOR_1_1_AND2_NUM160_OUT, XNOR_1_2_AND2_NUM160_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM160 (.ZN (XNOR_1_1_AND2_NUM160_OUT), .A1 (N154), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM160 (.ZN (XNOR_1_2_AND2_NUM160_OUT), .A1 (GND), .A2 (N528));
      NOR2_X1 XNOR_1_3_AND2_NUM160 (.ZN (N1020), .A1 (XNOR_1_1_AND2_NUM160_OUT), .A2 (XNOR_1_2_AND2_NUM160_OUT));
      wire XNOR_1_1_AND2_NUM161_OUT, XNOR_1_2_AND2_NUM161_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM161 (.ZN (XNOR_1_1_AND2_NUM161_OUT), .A1 (N171), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM161 (.ZN (XNOR_1_2_AND2_NUM161_OUT), .A1 (GND), .A2 (N273));
      NOR2_X1 XNOR_1_3_AND2_NUM161 (.ZN (N1023), .A1 (XNOR_1_1_AND2_NUM161_OUT), .A2 (XNOR_1_2_AND2_NUM161_OUT));
      wire XNOR_1_1_AND2_NUM162_OUT, XNOR_1_2_AND2_NUM162_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM162 (.ZN (XNOR_1_1_AND2_NUM162_OUT), .A1 (N171), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM162 (.ZN (XNOR_1_2_AND2_NUM162_OUT), .A1 (GND), .A2 (N290));
      NOR2_X1 XNOR_1_3_AND2_NUM162 (.ZN (N1026), .A1 (XNOR_1_1_AND2_NUM162_OUT), .A2 (XNOR_1_2_AND2_NUM162_OUT));
      wire XNOR_1_1_AND2_NUM163_OUT, XNOR_1_2_AND2_NUM163_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM163 (.ZN (XNOR_1_1_AND2_NUM163_OUT), .A1 (N171), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM163 (.ZN (XNOR_1_2_AND2_NUM163_OUT), .A1 (GND), .A2 (N307));
      NOR2_X1 XNOR_1_3_AND2_NUM163 (.ZN (N1029), .A1 (XNOR_1_1_AND2_NUM163_OUT), .A2 (XNOR_1_2_AND2_NUM163_OUT));
      wire XNOR_1_1_AND2_NUM164_OUT, XNOR_1_2_AND2_NUM164_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM164 (.ZN (XNOR_1_1_AND2_NUM164_OUT), .A1 (N171), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM164 (.ZN (XNOR_1_2_AND2_NUM164_OUT), .A1 (GND), .A2 (N324));
      NOR2_X1 XNOR_1_3_AND2_NUM164 (.ZN (N1032), .A1 (XNOR_1_1_AND2_NUM164_OUT), .A2 (XNOR_1_2_AND2_NUM164_OUT));
      wire XNOR_1_1_AND2_NUM165_OUT, XNOR_1_2_AND2_NUM165_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM165 (.ZN (XNOR_1_1_AND2_NUM165_OUT), .A1 (N171), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM165 (.ZN (XNOR_1_2_AND2_NUM165_OUT), .A1 (GND), .A2 (N341));
      NOR2_X1 XNOR_1_3_AND2_NUM165 (.ZN (N1035), .A1 (XNOR_1_1_AND2_NUM165_OUT), .A2 (XNOR_1_2_AND2_NUM165_OUT));
      wire XNOR_1_1_AND2_NUM166_OUT, XNOR_1_2_AND2_NUM166_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM166 (.ZN (XNOR_1_1_AND2_NUM166_OUT), .A1 (N171), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM166 (.ZN (XNOR_1_2_AND2_NUM166_OUT), .A1 (GND), .A2 (N358));
      NOR2_X1 XNOR_1_3_AND2_NUM166 (.ZN (N1038), .A1 (XNOR_1_1_AND2_NUM166_OUT), .A2 (XNOR_1_2_AND2_NUM166_OUT));
      wire XNOR_1_1_AND2_NUM167_OUT, XNOR_1_2_AND2_NUM167_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM167 (.ZN (XNOR_1_1_AND2_NUM167_OUT), .A1 (N171), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM167 (.ZN (XNOR_1_2_AND2_NUM167_OUT), .A1 (GND), .A2 (N375));
      NOR2_X1 XNOR_1_3_AND2_NUM167 (.ZN (N1041), .A1 (XNOR_1_1_AND2_NUM167_OUT), .A2 (XNOR_1_2_AND2_NUM167_OUT));
      wire XNOR_1_1_AND2_NUM168_OUT, XNOR_1_2_AND2_NUM168_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM168 (.ZN (XNOR_1_1_AND2_NUM168_OUT), .A1 (N171), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM168 (.ZN (XNOR_1_2_AND2_NUM168_OUT), .A1 (GND), .A2 (N392));
      NOR2_X1 XNOR_1_3_AND2_NUM168 (.ZN (N1044), .A1 (XNOR_1_1_AND2_NUM168_OUT), .A2 (XNOR_1_2_AND2_NUM168_OUT));
      wire XNOR_1_1_AND2_NUM169_OUT, XNOR_1_2_AND2_NUM169_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM169 (.ZN (XNOR_1_1_AND2_NUM169_OUT), .A1 (N171), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM169 (.ZN (XNOR_1_2_AND2_NUM169_OUT), .A1 (GND), .A2 (N409));
      NOR2_X1 XNOR_1_3_AND2_NUM169 (.ZN (N1047), .A1 (XNOR_1_1_AND2_NUM169_OUT), .A2 (XNOR_1_2_AND2_NUM169_OUT));
      wire XNOR_1_1_AND2_NUM170_OUT, XNOR_1_2_AND2_NUM170_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM170 (.ZN (XNOR_1_1_AND2_NUM170_OUT), .A1 (N171), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM170 (.ZN (XNOR_1_2_AND2_NUM170_OUT), .A1 (GND), .A2 (N426));
      NOR2_X1 XNOR_1_3_AND2_NUM170 (.ZN (N1050), .A1 (XNOR_1_1_AND2_NUM170_OUT), .A2 (XNOR_1_2_AND2_NUM170_OUT));
      wire XNOR_1_1_AND2_NUM171_OUT, XNOR_1_2_AND2_NUM171_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM171 (.ZN (XNOR_1_1_AND2_NUM171_OUT), .A1 (N171), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM171 (.ZN (XNOR_1_2_AND2_NUM171_OUT), .A1 (GND), .A2 (N443));
      NOR2_X1 XNOR_1_3_AND2_NUM171 (.ZN (N1053), .A1 (XNOR_1_1_AND2_NUM171_OUT), .A2 (XNOR_1_2_AND2_NUM171_OUT));
      wire XNOR_1_1_AND2_NUM172_OUT, XNOR_1_2_AND2_NUM172_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM172 (.ZN (XNOR_1_1_AND2_NUM172_OUT), .A1 (N171), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM172 (.ZN (XNOR_1_2_AND2_NUM172_OUT), .A1 (GND), .A2 (N460));
      NOR2_X1 XNOR_1_3_AND2_NUM172 (.ZN (N1056), .A1 (XNOR_1_1_AND2_NUM172_OUT), .A2 (XNOR_1_2_AND2_NUM172_OUT));
      wire XNOR_1_1_AND2_NUM173_OUT, XNOR_1_2_AND2_NUM173_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM173 (.ZN (XNOR_1_1_AND2_NUM173_OUT), .A1 (N171), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM173 (.ZN (XNOR_1_2_AND2_NUM173_OUT), .A1 (GND), .A2 (N477));
      NOR2_X1 XNOR_1_3_AND2_NUM173 (.ZN (N1059), .A1 (XNOR_1_1_AND2_NUM173_OUT), .A2 (XNOR_1_2_AND2_NUM173_OUT));
      wire XNOR_1_1_AND2_NUM174_OUT, XNOR_1_2_AND2_NUM174_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM174 (.ZN (XNOR_1_1_AND2_NUM174_OUT), .A1 (N171), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM174 (.ZN (XNOR_1_2_AND2_NUM174_OUT), .A1 (GND), .A2 (N494));
      NOR2_X1 XNOR_1_3_AND2_NUM174 (.ZN (N1062), .A1 (XNOR_1_1_AND2_NUM174_OUT), .A2 (XNOR_1_2_AND2_NUM174_OUT));
      wire XNOR_1_1_AND2_NUM175_OUT, XNOR_1_2_AND2_NUM175_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM175 (.ZN (XNOR_1_1_AND2_NUM175_OUT), .A1 (N171), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM175 (.ZN (XNOR_1_2_AND2_NUM175_OUT), .A1 (GND), .A2 (N511));
      NOR2_X1 XNOR_1_3_AND2_NUM175 (.ZN (N1065), .A1 (XNOR_1_1_AND2_NUM175_OUT), .A2 (XNOR_1_2_AND2_NUM175_OUT));
      wire XNOR_1_1_AND2_NUM176_OUT, XNOR_1_2_AND2_NUM176_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM176 (.ZN (XNOR_1_1_AND2_NUM176_OUT), .A1 (N171), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM176 (.ZN (XNOR_1_2_AND2_NUM176_OUT), .A1 (GND), .A2 (N528));
      NOR2_X1 XNOR_1_3_AND2_NUM176 (.ZN (N1068), .A1 (XNOR_1_1_AND2_NUM176_OUT), .A2 (XNOR_1_2_AND2_NUM176_OUT));
      wire XNOR_1_1_AND2_NUM177_OUT, XNOR_1_2_AND2_NUM177_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM177 (.ZN (XNOR_1_1_AND2_NUM177_OUT), .A1 (N188), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM177 (.ZN (XNOR_1_2_AND2_NUM177_OUT), .A1 (GND), .A2 (N273));
      NOR2_X1 XNOR_1_3_AND2_NUM177 (.ZN (N1071), .A1 (XNOR_1_1_AND2_NUM177_OUT), .A2 (XNOR_1_2_AND2_NUM177_OUT));
      wire XNOR_1_1_AND2_NUM178_OUT, XNOR_1_2_AND2_NUM178_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM178 (.ZN (XNOR_1_1_AND2_NUM178_OUT), .A1 (N188), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM178 (.ZN (XNOR_1_2_AND2_NUM178_OUT), .A1 (GND), .A2 (N290));
      NOR2_X1 XNOR_1_3_AND2_NUM178 (.ZN (N1074), .A1 (XNOR_1_1_AND2_NUM178_OUT), .A2 (XNOR_1_2_AND2_NUM178_OUT));
      wire XNOR_1_1_AND2_NUM179_OUT, XNOR_1_2_AND2_NUM179_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM179 (.ZN (XNOR_1_1_AND2_NUM179_OUT), .A1 (N188), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM179 (.ZN (XNOR_1_2_AND2_NUM179_OUT), .A1 (GND), .A2 (N307));
      NOR2_X1 XNOR_1_3_AND2_NUM179 (.ZN (N1077), .A1 (XNOR_1_1_AND2_NUM179_OUT), .A2 (XNOR_1_2_AND2_NUM179_OUT));
      wire XNOR_1_1_AND2_NUM180_OUT, XNOR_1_2_AND2_NUM180_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM180 (.ZN (XNOR_1_1_AND2_NUM180_OUT), .A1 (N188), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM180 (.ZN (XNOR_1_2_AND2_NUM180_OUT), .A1 (GND), .A2 (N324));
      NOR2_X1 XNOR_1_3_AND2_NUM180 (.ZN (N1080), .A1 (XNOR_1_1_AND2_NUM180_OUT), .A2 (XNOR_1_2_AND2_NUM180_OUT));
      wire XNOR_1_1_AND2_NUM181_OUT, XNOR_1_2_AND2_NUM181_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM181 (.ZN (XNOR_1_1_AND2_NUM181_OUT), .A1 (N188), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM181 (.ZN (XNOR_1_2_AND2_NUM181_OUT), .A1 (GND), .A2 (N341));
      NOR2_X1 XNOR_1_3_AND2_NUM181 (.ZN (N1083), .A1 (XNOR_1_1_AND2_NUM181_OUT), .A2 (XNOR_1_2_AND2_NUM181_OUT));
      wire XNOR_1_1_AND2_NUM182_OUT, XNOR_1_2_AND2_NUM182_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM182 (.ZN (XNOR_1_1_AND2_NUM182_OUT), .A1 (N188), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM182 (.ZN (XNOR_1_2_AND2_NUM182_OUT), .A1 (GND), .A2 (N358));
      NOR2_X1 XNOR_1_3_AND2_NUM182 (.ZN (N1086), .A1 (XNOR_1_1_AND2_NUM182_OUT), .A2 (XNOR_1_2_AND2_NUM182_OUT));
      wire XNOR_1_1_AND2_NUM183_OUT, XNOR_1_2_AND2_NUM183_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM183 (.ZN (XNOR_1_1_AND2_NUM183_OUT), .A1 (N188), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM183 (.ZN (XNOR_1_2_AND2_NUM183_OUT), .A1 (GND), .A2 (N375));
      NOR2_X1 XNOR_1_3_AND2_NUM183 (.ZN (N1089), .A1 (XNOR_1_1_AND2_NUM183_OUT), .A2 (XNOR_1_2_AND2_NUM183_OUT));
      wire XNOR_1_1_AND2_NUM184_OUT, XNOR_1_2_AND2_NUM184_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM184 (.ZN (XNOR_1_1_AND2_NUM184_OUT), .A1 (N188), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM184 (.ZN (XNOR_1_2_AND2_NUM184_OUT), .A1 (GND), .A2 (N392));
      NOR2_X1 XNOR_1_3_AND2_NUM184 (.ZN (N1092), .A1 (XNOR_1_1_AND2_NUM184_OUT), .A2 (XNOR_1_2_AND2_NUM184_OUT));
      wire XNOR_1_1_AND2_NUM185_OUT, XNOR_1_2_AND2_NUM185_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM185 (.ZN (XNOR_1_1_AND2_NUM185_OUT), .A1 (N188), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM185 (.ZN (XNOR_1_2_AND2_NUM185_OUT), .A1 (GND), .A2 (N409));
      NOR2_X1 XNOR_1_3_AND2_NUM185 (.ZN (N1095), .A1 (XNOR_1_1_AND2_NUM185_OUT), .A2 (XNOR_1_2_AND2_NUM185_OUT));
      wire XNOR_1_1_AND2_NUM186_OUT, XNOR_1_2_AND2_NUM186_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM186 (.ZN (XNOR_1_1_AND2_NUM186_OUT), .A1 (N188), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM186 (.ZN (XNOR_1_2_AND2_NUM186_OUT), .A1 (GND), .A2 (N426));
      NOR2_X1 XNOR_1_3_AND2_NUM186 (.ZN (N1098), .A1 (XNOR_1_1_AND2_NUM186_OUT), .A2 (XNOR_1_2_AND2_NUM186_OUT));
      wire XNOR_1_1_AND2_NUM187_OUT, XNOR_1_2_AND2_NUM187_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM187 (.ZN (XNOR_1_1_AND2_NUM187_OUT), .A1 (N188), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM187 (.ZN (XNOR_1_2_AND2_NUM187_OUT), .A1 (GND), .A2 (N443));
      NOR2_X1 XNOR_1_3_AND2_NUM187 (.ZN (N1101), .A1 (XNOR_1_1_AND2_NUM187_OUT), .A2 (XNOR_1_2_AND2_NUM187_OUT));
      wire XNOR_1_1_AND2_NUM188_OUT, XNOR_1_2_AND2_NUM188_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM188 (.ZN (XNOR_1_1_AND2_NUM188_OUT), .A1 (N188), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM188 (.ZN (XNOR_1_2_AND2_NUM188_OUT), .A1 (GND), .A2 (N460));
      NOR2_X1 XNOR_1_3_AND2_NUM188 (.ZN (N1104), .A1 (XNOR_1_1_AND2_NUM188_OUT), .A2 (XNOR_1_2_AND2_NUM188_OUT));
      wire XNOR_1_1_AND2_NUM189_OUT, XNOR_1_2_AND2_NUM189_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM189 (.ZN (XNOR_1_1_AND2_NUM189_OUT), .A1 (N188), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM189 (.ZN (XNOR_1_2_AND2_NUM189_OUT), .A1 (GND), .A2 (N477));
      NOR2_X1 XNOR_1_3_AND2_NUM189 (.ZN (N1107), .A1 (XNOR_1_1_AND2_NUM189_OUT), .A2 (XNOR_1_2_AND2_NUM189_OUT));
      wire XNOR_1_1_AND2_NUM190_OUT, XNOR_1_2_AND2_NUM190_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM190 (.ZN (XNOR_1_1_AND2_NUM190_OUT), .A1 (N188), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM190 (.ZN (XNOR_1_2_AND2_NUM190_OUT), .A1 (GND), .A2 (N494));
      NOR2_X1 XNOR_1_3_AND2_NUM190 (.ZN (N1110), .A1 (XNOR_1_1_AND2_NUM190_OUT), .A2 (XNOR_1_2_AND2_NUM190_OUT));
      wire XNOR_1_1_AND2_NUM191_OUT, XNOR_1_2_AND2_NUM191_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM191 (.ZN (XNOR_1_1_AND2_NUM191_OUT), .A1 (N188), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM191 (.ZN (XNOR_1_2_AND2_NUM191_OUT), .A1 (GND), .A2 (N511));
      NOR2_X1 XNOR_1_3_AND2_NUM191 (.ZN (N1113), .A1 (XNOR_1_1_AND2_NUM191_OUT), .A2 (XNOR_1_2_AND2_NUM191_OUT));
      wire XNOR_1_1_AND2_NUM192_OUT, XNOR_1_2_AND2_NUM192_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM192 (.ZN (XNOR_1_1_AND2_NUM192_OUT), .A1 (N188), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM192 (.ZN (XNOR_1_2_AND2_NUM192_OUT), .A1 (GND), .A2 (N528));
      NOR2_X1 XNOR_1_3_AND2_NUM192 (.ZN (N1116), .A1 (XNOR_1_1_AND2_NUM192_OUT), .A2 (XNOR_1_2_AND2_NUM192_OUT));
      wire XNOR_1_1_AND2_NUM193_OUT, XNOR_1_2_AND2_NUM193_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM193 (.ZN (XNOR_1_1_AND2_NUM193_OUT), .A1 (N205), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM193 (.ZN (XNOR_1_2_AND2_NUM193_OUT), .A1 (GND), .A2 (N273));
      NOR2_X1 XNOR_1_3_AND2_NUM193 (.ZN (N1119), .A1 (XNOR_1_1_AND2_NUM193_OUT), .A2 (XNOR_1_2_AND2_NUM193_OUT));
      wire XNOR_1_1_AND2_NUM194_OUT, XNOR_1_2_AND2_NUM194_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM194 (.ZN (XNOR_1_1_AND2_NUM194_OUT), .A1 (N205), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM194 (.ZN (XNOR_1_2_AND2_NUM194_OUT), .A1 (GND), .A2 (N290));
      NOR2_X1 XNOR_1_3_AND2_NUM194 (.ZN (N1122), .A1 (XNOR_1_1_AND2_NUM194_OUT), .A2 (XNOR_1_2_AND2_NUM194_OUT));
      wire XNOR_1_1_AND2_NUM195_OUT, XNOR_1_2_AND2_NUM195_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM195 (.ZN (XNOR_1_1_AND2_NUM195_OUT), .A1 (N205), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM195 (.ZN (XNOR_1_2_AND2_NUM195_OUT), .A1 (GND), .A2 (N307));
      NOR2_X1 XNOR_1_3_AND2_NUM195 (.ZN (N1125), .A1 (XNOR_1_1_AND2_NUM195_OUT), .A2 (XNOR_1_2_AND2_NUM195_OUT));
      wire XNOR_1_1_AND2_NUM196_OUT, XNOR_1_2_AND2_NUM196_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM196 (.ZN (XNOR_1_1_AND2_NUM196_OUT), .A1 (N205), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM196 (.ZN (XNOR_1_2_AND2_NUM196_OUT), .A1 (GND), .A2 (N324));
      NOR2_X1 XNOR_1_3_AND2_NUM196 (.ZN (N1128), .A1 (XNOR_1_1_AND2_NUM196_OUT), .A2 (XNOR_1_2_AND2_NUM196_OUT));
      wire XNOR_1_1_AND2_NUM197_OUT, XNOR_1_2_AND2_NUM197_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM197 (.ZN (XNOR_1_1_AND2_NUM197_OUT), .A1 (N205), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM197 (.ZN (XNOR_1_2_AND2_NUM197_OUT), .A1 (GND), .A2 (N341));
      NOR2_X1 XNOR_1_3_AND2_NUM197 (.ZN (N1131), .A1 (XNOR_1_1_AND2_NUM197_OUT), .A2 (XNOR_1_2_AND2_NUM197_OUT));
      wire XNOR_1_1_AND2_NUM198_OUT, XNOR_1_2_AND2_NUM198_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM198 (.ZN (XNOR_1_1_AND2_NUM198_OUT), .A1 (N205), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM198 (.ZN (XNOR_1_2_AND2_NUM198_OUT), .A1 (GND), .A2 (N358));
      NOR2_X1 XNOR_1_3_AND2_NUM198 (.ZN (N1134), .A1 (XNOR_1_1_AND2_NUM198_OUT), .A2 (XNOR_1_2_AND2_NUM198_OUT));
      wire XNOR_1_1_AND2_NUM199_OUT, XNOR_1_2_AND2_NUM199_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM199 (.ZN (XNOR_1_1_AND2_NUM199_OUT), .A1 (N205), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM199 (.ZN (XNOR_1_2_AND2_NUM199_OUT), .A1 (GND), .A2 (N375));
      NOR2_X1 XNOR_1_3_AND2_NUM199 (.ZN (N1137), .A1 (XNOR_1_1_AND2_NUM199_OUT), .A2 (XNOR_1_2_AND2_NUM199_OUT));
      wire XNOR_1_1_AND2_NUM200_OUT, XNOR_1_2_AND2_NUM200_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM200 (.ZN (XNOR_1_1_AND2_NUM200_OUT), .A1 (N205), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM200 (.ZN (XNOR_1_2_AND2_NUM200_OUT), .A1 (GND), .A2 (N392));
      NOR2_X1 XNOR_1_3_AND2_NUM200 (.ZN (N1140), .A1 (XNOR_1_1_AND2_NUM200_OUT), .A2 (XNOR_1_2_AND2_NUM200_OUT));
      wire XNOR_1_1_AND2_NUM201_OUT, XNOR_1_2_AND2_NUM201_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM201 (.ZN (XNOR_1_1_AND2_NUM201_OUT), .A1 (N205), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM201 (.ZN (XNOR_1_2_AND2_NUM201_OUT), .A1 (GND), .A2 (N409));
      NOR2_X1 XNOR_1_3_AND2_NUM201 (.ZN (N1143), .A1 (XNOR_1_1_AND2_NUM201_OUT), .A2 (XNOR_1_2_AND2_NUM201_OUT));
      wire XNOR_1_1_AND2_NUM202_OUT, XNOR_1_2_AND2_NUM202_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM202 (.ZN (XNOR_1_1_AND2_NUM202_OUT), .A1 (N205), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM202 (.ZN (XNOR_1_2_AND2_NUM202_OUT), .A1 (GND), .A2 (N426));
      NOR2_X1 XNOR_1_3_AND2_NUM202 (.ZN (N1146), .A1 (XNOR_1_1_AND2_NUM202_OUT), .A2 (XNOR_1_2_AND2_NUM202_OUT));
      wire XNOR_1_1_AND2_NUM203_OUT, XNOR_1_2_AND2_NUM203_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM203 (.ZN (XNOR_1_1_AND2_NUM203_OUT), .A1 (N205), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM203 (.ZN (XNOR_1_2_AND2_NUM203_OUT), .A1 (GND), .A2 (N443));
      NOR2_X1 XNOR_1_3_AND2_NUM203 (.ZN (N1149), .A1 (XNOR_1_1_AND2_NUM203_OUT), .A2 (XNOR_1_2_AND2_NUM203_OUT));
      wire XNOR_1_1_AND2_NUM204_OUT, XNOR_1_2_AND2_NUM204_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM204 (.ZN (XNOR_1_1_AND2_NUM204_OUT), .A1 (N205), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM204 (.ZN (XNOR_1_2_AND2_NUM204_OUT), .A1 (GND), .A2 (N460));
      NOR2_X1 XNOR_1_3_AND2_NUM204 (.ZN (N1152), .A1 (XNOR_1_1_AND2_NUM204_OUT), .A2 (XNOR_1_2_AND2_NUM204_OUT));
      wire XNOR_1_1_AND2_NUM205_OUT, XNOR_1_2_AND2_NUM205_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM205 (.ZN (XNOR_1_1_AND2_NUM205_OUT), .A1 (N205), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM205 (.ZN (XNOR_1_2_AND2_NUM205_OUT), .A1 (GND), .A2 (N477));
      NOR2_X1 XNOR_1_3_AND2_NUM205 (.ZN (N1155), .A1 (XNOR_1_1_AND2_NUM205_OUT), .A2 (XNOR_1_2_AND2_NUM205_OUT));
      wire XNOR_1_1_AND2_NUM206_OUT, XNOR_1_2_AND2_NUM206_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM206 (.ZN (XNOR_1_1_AND2_NUM206_OUT), .A1 (N205), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM206 (.ZN (XNOR_1_2_AND2_NUM206_OUT), .A1 (GND), .A2 (N494));
      NOR2_X1 XNOR_1_3_AND2_NUM206 (.ZN (N1158), .A1 (XNOR_1_1_AND2_NUM206_OUT), .A2 (XNOR_1_2_AND2_NUM206_OUT));
      wire XNOR_1_1_AND2_NUM207_OUT, XNOR_1_2_AND2_NUM207_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM207 (.ZN (XNOR_1_1_AND2_NUM207_OUT), .A1 (N205), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM207 (.ZN (XNOR_1_2_AND2_NUM207_OUT), .A1 (GND), .A2 (N511));
      NOR2_X1 XNOR_1_3_AND2_NUM207 (.ZN (N1161), .A1 (XNOR_1_1_AND2_NUM207_OUT), .A2 (XNOR_1_2_AND2_NUM207_OUT));
      wire XNOR_1_1_AND2_NUM208_OUT, XNOR_1_2_AND2_NUM208_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM208 (.ZN (XNOR_1_1_AND2_NUM208_OUT), .A1 (N205), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM208 (.ZN (XNOR_1_2_AND2_NUM208_OUT), .A1 (GND), .A2 (N528));
      NOR2_X1 XNOR_1_3_AND2_NUM208 (.ZN (N1164), .A1 (XNOR_1_1_AND2_NUM208_OUT), .A2 (XNOR_1_2_AND2_NUM208_OUT));
      wire XNOR_1_1_AND2_NUM209_OUT, XNOR_1_2_AND2_NUM209_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM209 (.ZN (XNOR_1_1_AND2_NUM209_OUT), .A1 (N222), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM209 (.ZN (XNOR_1_2_AND2_NUM209_OUT), .A1 (GND), .A2 (N273));
      NOR2_X1 XNOR_1_3_AND2_NUM209 (.ZN (N1167), .A1 (XNOR_1_1_AND2_NUM209_OUT), .A2 (XNOR_1_2_AND2_NUM209_OUT));
      wire XNOR_1_1_AND2_NUM210_OUT, XNOR_1_2_AND2_NUM210_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM210 (.ZN (XNOR_1_1_AND2_NUM210_OUT), .A1 (N222), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM210 (.ZN (XNOR_1_2_AND2_NUM210_OUT), .A1 (GND), .A2 (N290));
      NOR2_X1 XNOR_1_3_AND2_NUM210 (.ZN (N1170), .A1 (XNOR_1_1_AND2_NUM210_OUT), .A2 (XNOR_1_2_AND2_NUM210_OUT));
      wire XNOR_1_1_AND2_NUM211_OUT, XNOR_1_2_AND2_NUM211_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM211 (.ZN (XNOR_1_1_AND2_NUM211_OUT), .A1 (N222), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM211 (.ZN (XNOR_1_2_AND2_NUM211_OUT), .A1 (GND), .A2 (N307));
      NOR2_X1 XNOR_1_3_AND2_NUM211 (.ZN (N1173), .A1 (XNOR_1_1_AND2_NUM211_OUT), .A2 (XNOR_1_2_AND2_NUM211_OUT));
      wire XNOR_1_1_AND2_NUM212_OUT, XNOR_1_2_AND2_NUM212_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM212 (.ZN (XNOR_1_1_AND2_NUM212_OUT), .A1 (N222), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM212 (.ZN (XNOR_1_2_AND2_NUM212_OUT), .A1 (GND), .A2 (N324));
      NOR2_X1 XNOR_1_3_AND2_NUM212 (.ZN (N1176), .A1 (XNOR_1_1_AND2_NUM212_OUT), .A2 (XNOR_1_2_AND2_NUM212_OUT));
      wire XNOR_1_1_AND2_NUM213_OUT, XNOR_1_2_AND2_NUM213_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM213 (.ZN (XNOR_1_1_AND2_NUM213_OUT), .A1 (N222), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM213 (.ZN (XNOR_1_2_AND2_NUM213_OUT), .A1 (GND), .A2 (N341));
      NOR2_X1 XNOR_1_3_AND2_NUM213 (.ZN (N1179), .A1 (XNOR_1_1_AND2_NUM213_OUT), .A2 (XNOR_1_2_AND2_NUM213_OUT));
      wire XNOR_1_1_AND2_NUM214_OUT, XNOR_1_2_AND2_NUM214_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM214 (.ZN (XNOR_1_1_AND2_NUM214_OUT), .A1 (N222), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM214 (.ZN (XNOR_1_2_AND2_NUM214_OUT), .A1 (GND), .A2 (N358));
      NOR2_X1 XNOR_1_3_AND2_NUM214 (.ZN (N1182), .A1 (XNOR_1_1_AND2_NUM214_OUT), .A2 (XNOR_1_2_AND2_NUM214_OUT));
      wire XNOR_1_1_AND2_NUM215_OUT, XNOR_1_2_AND2_NUM215_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM215 (.ZN (XNOR_1_1_AND2_NUM215_OUT), .A1 (N222), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM215 (.ZN (XNOR_1_2_AND2_NUM215_OUT), .A1 (GND), .A2 (N375));
      NOR2_X1 XNOR_1_3_AND2_NUM215 (.ZN (N1185), .A1 (XNOR_1_1_AND2_NUM215_OUT), .A2 (XNOR_1_2_AND2_NUM215_OUT));
      wire XNOR_1_1_AND2_NUM216_OUT, XNOR_1_2_AND2_NUM216_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM216 (.ZN (XNOR_1_1_AND2_NUM216_OUT), .A1 (N222), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM216 (.ZN (XNOR_1_2_AND2_NUM216_OUT), .A1 (GND), .A2 (N392));
      NOR2_X1 XNOR_1_3_AND2_NUM216 (.ZN (N1188), .A1 (XNOR_1_1_AND2_NUM216_OUT), .A2 (XNOR_1_2_AND2_NUM216_OUT));
      wire XNOR_1_1_AND2_NUM217_OUT, XNOR_1_2_AND2_NUM217_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM217 (.ZN (XNOR_1_1_AND2_NUM217_OUT), .A1 (N222), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM217 (.ZN (XNOR_1_2_AND2_NUM217_OUT), .A1 (GND), .A2 (N409));
      NOR2_X1 XNOR_1_3_AND2_NUM217 (.ZN (N1191), .A1 (XNOR_1_1_AND2_NUM217_OUT), .A2 (XNOR_1_2_AND2_NUM217_OUT));
      wire XNOR_1_1_AND2_NUM218_OUT, XNOR_1_2_AND2_NUM218_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM218 (.ZN (XNOR_1_1_AND2_NUM218_OUT), .A1 (N222), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM218 (.ZN (XNOR_1_2_AND2_NUM218_OUT), .A1 (GND), .A2 (N426));
      NOR2_X1 XNOR_1_3_AND2_NUM218 (.ZN (N1194), .A1 (XNOR_1_1_AND2_NUM218_OUT), .A2 (XNOR_1_2_AND2_NUM218_OUT));
      wire XNOR_1_1_AND2_NUM219_OUT, XNOR_1_2_AND2_NUM219_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM219 (.ZN (XNOR_1_1_AND2_NUM219_OUT), .A1 (N222), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM219 (.ZN (XNOR_1_2_AND2_NUM219_OUT), .A1 (GND), .A2 (N443));
      NOR2_X1 XNOR_1_3_AND2_NUM219 (.ZN (N1197), .A1 (XNOR_1_1_AND2_NUM219_OUT), .A2 (XNOR_1_2_AND2_NUM219_OUT));
      wire XNOR_1_1_AND2_NUM220_OUT, XNOR_1_2_AND2_NUM220_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM220 (.ZN (XNOR_1_1_AND2_NUM220_OUT), .A1 (N222), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM220 (.ZN (XNOR_1_2_AND2_NUM220_OUT), .A1 (GND), .A2 (N460));
      NOR2_X1 XNOR_1_3_AND2_NUM220 (.ZN (N1200), .A1 (XNOR_1_1_AND2_NUM220_OUT), .A2 (XNOR_1_2_AND2_NUM220_OUT));
      wire XNOR_1_1_AND2_NUM221_OUT, XNOR_1_2_AND2_NUM221_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM221 (.ZN (XNOR_1_1_AND2_NUM221_OUT), .A1 (N222), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM221 (.ZN (XNOR_1_2_AND2_NUM221_OUT), .A1 (GND), .A2 (N477));
      NOR2_X1 XNOR_1_3_AND2_NUM221 (.ZN (N1203), .A1 (XNOR_1_1_AND2_NUM221_OUT), .A2 (XNOR_1_2_AND2_NUM221_OUT));
      wire XNOR_1_1_AND2_NUM222_OUT, XNOR_1_2_AND2_NUM222_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM222 (.ZN (XNOR_1_1_AND2_NUM222_OUT), .A1 (N222), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM222 (.ZN (XNOR_1_2_AND2_NUM222_OUT), .A1 (GND), .A2 (N494));
      NOR2_X1 XNOR_1_3_AND2_NUM222 (.ZN (N1206), .A1 (XNOR_1_1_AND2_NUM222_OUT), .A2 (XNOR_1_2_AND2_NUM222_OUT));
      wire XNOR_1_1_AND2_NUM223_OUT, XNOR_1_2_AND2_NUM223_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM223 (.ZN (XNOR_1_1_AND2_NUM223_OUT), .A1 (N222), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM223 (.ZN (XNOR_1_2_AND2_NUM223_OUT), .A1 (GND), .A2 (N511));
      NOR2_X1 XNOR_1_3_AND2_NUM223 (.ZN (N1209), .A1 (XNOR_1_1_AND2_NUM223_OUT), .A2 (XNOR_1_2_AND2_NUM223_OUT));
      wire XNOR_1_1_AND2_NUM224_OUT, XNOR_1_2_AND2_NUM224_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM224 (.ZN (XNOR_1_1_AND2_NUM224_OUT), .A1 (N222), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM224 (.ZN (XNOR_1_2_AND2_NUM224_OUT), .A1 (GND), .A2 (N528));
      NOR2_X1 XNOR_1_3_AND2_NUM224 (.ZN (N1212), .A1 (XNOR_1_1_AND2_NUM224_OUT), .A2 (XNOR_1_2_AND2_NUM224_OUT));
      wire XNOR_1_1_AND2_NUM225_OUT, XNOR_1_2_AND2_NUM225_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM225 (.ZN (XNOR_1_1_AND2_NUM225_OUT), .A1 (N239), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM225 (.ZN (XNOR_1_2_AND2_NUM225_OUT), .A1 (GND), .A2 (N273));
      NOR2_X1 XNOR_1_3_AND2_NUM225 (.ZN (N1215), .A1 (XNOR_1_1_AND2_NUM225_OUT), .A2 (XNOR_1_2_AND2_NUM225_OUT));
      wire XNOR_1_1_AND2_NUM226_OUT, XNOR_1_2_AND2_NUM226_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM226 (.ZN (XNOR_1_1_AND2_NUM226_OUT), .A1 (N239), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM226 (.ZN (XNOR_1_2_AND2_NUM226_OUT), .A1 (GND), .A2 (N290));
      NOR2_X1 XNOR_1_3_AND2_NUM226 (.ZN (N1218), .A1 (XNOR_1_1_AND2_NUM226_OUT), .A2 (XNOR_1_2_AND2_NUM226_OUT));
      wire XNOR_1_1_AND2_NUM227_OUT, XNOR_1_2_AND2_NUM227_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM227 (.ZN (XNOR_1_1_AND2_NUM227_OUT), .A1 (N239), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM227 (.ZN (XNOR_1_2_AND2_NUM227_OUT), .A1 (GND), .A2 (N307));
      NOR2_X1 XNOR_1_3_AND2_NUM227 (.ZN (N1221), .A1 (XNOR_1_1_AND2_NUM227_OUT), .A2 (XNOR_1_2_AND2_NUM227_OUT));
      wire XNOR_1_1_AND2_NUM228_OUT, XNOR_1_2_AND2_NUM228_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM228 (.ZN (XNOR_1_1_AND2_NUM228_OUT), .A1 (N239), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM228 (.ZN (XNOR_1_2_AND2_NUM228_OUT), .A1 (GND), .A2 (N324));
      NOR2_X1 XNOR_1_3_AND2_NUM228 (.ZN (N1224), .A1 (XNOR_1_1_AND2_NUM228_OUT), .A2 (XNOR_1_2_AND2_NUM228_OUT));
      wire XNOR_1_1_AND2_NUM229_OUT, XNOR_1_2_AND2_NUM229_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM229 (.ZN (XNOR_1_1_AND2_NUM229_OUT), .A1 (N239), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM229 (.ZN (XNOR_1_2_AND2_NUM229_OUT), .A1 (GND), .A2 (N341));
      NOR2_X1 XNOR_1_3_AND2_NUM229 (.ZN (N1227), .A1 (XNOR_1_1_AND2_NUM229_OUT), .A2 (XNOR_1_2_AND2_NUM229_OUT));
      wire XNOR_1_1_AND2_NUM230_OUT, XNOR_1_2_AND2_NUM230_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM230 (.ZN (XNOR_1_1_AND2_NUM230_OUT), .A1 (N239), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM230 (.ZN (XNOR_1_2_AND2_NUM230_OUT), .A1 (GND), .A2 (N358));
      NOR2_X1 XNOR_1_3_AND2_NUM230 (.ZN (N1230), .A1 (XNOR_1_1_AND2_NUM230_OUT), .A2 (XNOR_1_2_AND2_NUM230_OUT));
      wire XNOR_1_1_AND2_NUM231_OUT, XNOR_1_2_AND2_NUM231_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM231 (.ZN (XNOR_1_1_AND2_NUM231_OUT), .A1 (N239), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM231 (.ZN (XNOR_1_2_AND2_NUM231_OUT), .A1 (GND), .A2 (N375));
      NOR2_X1 XNOR_1_3_AND2_NUM231 (.ZN (N1233), .A1 (XNOR_1_1_AND2_NUM231_OUT), .A2 (XNOR_1_2_AND2_NUM231_OUT));
      wire XNOR_1_1_AND2_NUM232_OUT, XNOR_1_2_AND2_NUM232_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM232 (.ZN (XNOR_1_1_AND2_NUM232_OUT), .A1 (N239), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM232 (.ZN (XNOR_1_2_AND2_NUM232_OUT), .A1 (GND), .A2 (N392));
      NOR2_X1 XNOR_1_3_AND2_NUM232 (.ZN (N1236), .A1 (XNOR_1_1_AND2_NUM232_OUT), .A2 (XNOR_1_2_AND2_NUM232_OUT));
      wire XNOR_1_1_AND2_NUM233_OUT, XNOR_1_2_AND2_NUM233_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM233 (.ZN (XNOR_1_1_AND2_NUM233_OUT), .A1 (N239), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM233 (.ZN (XNOR_1_2_AND2_NUM233_OUT), .A1 (GND), .A2 (N409));
      NOR2_X1 XNOR_1_3_AND2_NUM233 (.ZN (N1239), .A1 (XNOR_1_1_AND2_NUM233_OUT), .A2 (XNOR_1_2_AND2_NUM233_OUT));
      wire XNOR_1_1_AND2_NUM234_OUT, XNOR_1_2_AND2_NUM234_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM234 (.ZN (XNOR_1_1_AND2_NUM234_OUT), .A1 (N239), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM234 (.ZN (XNOR_1_2_AND2_NUM234_OUT), .A1 (GND), .A2 (N426));
      NOR2_X1 XNOR_1_3_AND2_NUM234 (.ZN (N1242), .A1 (XNOR_1_1_AND2_NUM234_OUT), .A2 (XNOR_1_2_AND2_NUM234_OUT));
      wire XNOR_1_1_AND2_NUM235_OUT, XNOR_1_2_AND2_NUM235_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM235 (.ZN (XNOR_1_1_AND2_NUM235_OUT), .A1 (N239), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM235 (.ZN (XNOR_1_2_AND2_NUM235_OUT), .A1 (GND), .A2 (N443));
      NOR2_X1 XNOR_1_3_AND2_NUM235 (.ZN (N1245), .A1 (XNOR_1_1_AND2_NUM235_OUT), .A2 (XNOR_1_2_AND2_NUM235_OUT));
      wire XNOR_1_1_AND2_NUM236_OUT, XNOR_1_2_AND2_NUM236_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM236 (.ZN (XNOR_1_1_AND2_NUM236_OUT), .A1 (N239), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM236 (.ZN (XNOR_1_2_AND2_NUM236_OUT), .A1 (GND), .A2 (N460));
      NOR2_X1 XNOR_1_3_AND2_NUM236 (.ZN (N1248), .A1 (XNOR_1_1_AND2_NUM236_OUT), .A2 (XNOR_1_2_AND2_NUM236_OUT));
      wire XNOR_1_1_AND2_NUM237_OUT, XNOR_1_2_AND2_NUM237_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM237 (.ZN (XNOR_1_1_AND2_NUM237_OUT), .A1 (N239), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM237 (.ZN (XNOR_1_2_AND2_NUM237_OUT), .A1 (GND), .A2 (N477));
      NOR2_X1 XNOR_1_3_AND2_NUM237 (.ZN (N1251), .A1 (XNOR_1_1_AND2_NUM237_OUT), .A2 (XNOR_1_2_AND2_NUM237_OUT));
      wire XNOR_1_1_AND2_NUM238_OUT, XNOR_1_2_AND2_NUM238_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM238 (.ZN (XNOR_1_1_AND2_NUM238_OUT), .A1 (N239), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM238 (.ZN (XNOR_1_2_AND2_NUM238_OUT), .A1 (GND), .A2 (N494));
      NOR2_X1 XNOR_1_3_AND2_NUM238 (.ZN (N1254), .A1 (XNOR_1_1_AND2_NUM238_OUT), .A2 (XNOR_1_2_AND2_NUM238_OUT));
      wire XNOR_1_1_AND2_NUM239_OUT, XNOR_1_2_AND2_NUM239_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM239 (.ZN (XNOR_1_1_AND2_NUM239_OUT), .A1 (N239), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM239 (.ZN (XNOR_1_2_AND2_NUM239_OUT), .A1 (GND), .A2 (N511));
      NOR2_X1 XNOR_1_3_AND2_NUM239 (.ZN (N1257), .A1 (XNOR_1_1_AND2_NUM239_OUT), .A2 (XNOR_1_2_AND2_NUM239_OUT));
      wire XNOR_1_1_AND2_NUM240_OUT, XNOR_1_2_AND2_NUM240_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM240 (.ZN (XNOR_1_1_AND2_NUM240_OUT), .A1 (N239), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM240 (.ZN (XNOR_1_2_AND2_NUM240_OUT), .A1 (GND), .A2 (N528));
      NOR2_X1 XNOR_1_3_AND2_NUM240 (.ZN (N1260), .A1 (XNOR_1_1_AND2_NUM240_OUT), .A2 (XNOR_1_2_AND2_NUM240_OUT));
      wire XNOR_1_1_AND2_NUM241_OUT, XNOR_1_2_AND2_NUM241_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM241 (.ZN (XNOR_1_1_AND2_NUM241_OUT), .A1 (N256), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM241 (.ZN (XNOR_1_2_AND2_NUM241_OUT), .A1 (GND), .A2 (N273));
      NOR2_X1 XNOR_1_3_AND2_NUM241 (.ZN (N1263), .A1 (XNOR_1_1_AND2_NUM241_OUT), .A2 (XNOR_1_2_AND2_NUM241_OUT));
      wire XNOR_1_1_AND2_NUM242_OUT, XNOR_1_2_AND2_NUM242_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM242 (.ZN (XNOR_1_1_AND2_NUM242_OUT), .A1 (N256), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM242 (.ZN (XNOR_1_2_AND2_NUM242_OUT), .A1 (GND), .A2 (N290));
      NOR2_X1 XNOR_1_3_AND2_NUM242 (.ZN (N1266), .A1 (XNOR_1_1_AND2_NUM242_OUT), .A2 (XNOR_1_2_AND2_NUM242_OUT));
      wire XNOR_1_1_AND2_NUM243_OUT, XNOR_1_2_AND2_NUM243_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM243 (.ZN (XNOR_1_1_AND2_NUM243_OUT), .A1 (N256), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM243 (.ZN (XNOR_1_2_AND2_NUM243_OUT), .A1 (GND), .A2 (N307));
      NOR2_X1 XNOR_1_3_AND2_NUM243 (.ZN (N1269), .A1 (XNOR_1_1_AND2_NUM243_OUT), .A2 (XNOR_1_2_AND2_NUM243_OUT));
      wire XNOR_1_1_AND2_NUM244_OUT, XNOR_1_2_AND2_NUM244_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM244 (.ZN (XNOR_1_1_AND2_NUM244_OUT), .A1 (N256), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM244 (.ZN (XNOR_1_2_AND2_NUM244_OUT), .A1 (GND), .A2 (N324));
      NOR2_X1 XNOR_1_3_AND2_NUM244 (.ZN (N1272), .A1 (XNOR_1_1_AND2_NUM244_OUT), .A2 (XNOR_1_2_AND2_NUM244_OUT));
      wire XNOR_1_1_AND2_NUM245_OUT, XNOR_1_2_AND2_NUM245_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM245 (.ZN (XNOR_1_1_AND2_NUM245_OUT), .A1 (N256), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM245 (.ZN (XNOR_1_2_AND2_NUM245_OUT), .A1 (GND), .A2 (N341));
      NOR2_X1 XNOR_1_3_AND2_NUM245 (.ZN (N1275), .A1 (XNOR_1_1_AND2_NUM245_OUT), .A2 (XNOR_1_2_AND2_NUM245_OUT));
      wire XNOR_1_1_AND2_NUM246_OUT, XNOR_1_2_AND2_NUM246_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM246 (.ZN (XNOR_1_1_AND2_NUM246_OUT), .A1 (N256), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM246 (.ZN (XNOR_1_2_AND2_NUM246_OUT), .A1 (GND), .A2 (N358));
      NOR2_X1 XNOR_1_3_AND2_NUM246 (.ZN (N1278), .A1 (XNOR_1_1_AND2_NUM246_OUT), .A2 (XNOR_1_2_AND2_NUM246_OUT));
      wire XNOR_1_1_AND2_NUM247_OUT, XNOR_1_2_AND2_NUM247_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM247 (.ZN (XNOR_1_1_AND2_NUM247_OUT), .A1 (N256), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM247 (.ZN (XNOR_1_2_AND2_NUM247_OUT), .A1 (GND), .A2 (N375));
      NOR2_X1 XNOR_1_3_AND2_NUM247 (.ZN (N1281), .A1 (XNOR_1_1_AND2_NUM247_OUT), .A2 (XNOR_1_2_AND2_NUM247_OUT));
      wire XNOR_1_1_AND2_NUM248_OUT, XNOR_1_2_AND2_NUM248_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM248 (.ZN (XNOR_1_1_AND2_NUM248_OUT), .A1 (N256), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM248 (.ZN (XNOR_1_2_AND2_NUM248_OUT), .A1 (GND), .A2 (N392));
      NOR2_X1 XNOR_1_3_AND2_NUM248 (.ZN (N1284), .A1 (XNOR_1_1_AND2_NUM248_OUT), .A2 (XNOR_1_2_AND2_NUM248_OUT));
      wire XNOR_1_1_AND2_NUM249_OUT, XNOR_1_2_AND2_NUM249_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM249 (.ZN (XNOR_1_1_AND2_NUM249_OUT), .A1 (N256), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM249 (.ZN (XNOR_1_2_AND2_NUM249_OUT), .A1 (GND), .A2 (N409));
      NOR2_X1 XNOR_1_3_AND2_NUM249 (.ZN (N1287), .A1 (XNOR_1_1_AND2_NUM249_OUT), .A2 (XNOR_1_2_AND2_NUM249_OUT));
      wire XNOR_1_1_AND2_NUM250_OUT, XNOR_1_2_AND2_NUM250_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM250 (.ZN (XNOR_1_1_AND2_NUM250_OUT), .A1 (N256), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM250 (.ZN (XNOR_1_2_AND2_NUM250_OUT), .A1 (GND), .A2 (N426));
      NOR2_X1 XNOR_1_3_AND2_NUM250 (.ZN (N1290), .A1 (XNOR_1_1_AND2_NUM250_OUT), .A2 (XNOR_1_2_AND2_NUM250_OUT));
      wire XNOR_1_1_AND2_NUM251_OUT, XNOR_1_2_AND2_NUM251_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM251 (.ZN (XNOR_1_1_AND2_NUM251_OUT), .A1 (N256), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM251 (.ZN (XNOR_1_2_AND2_NUM251_OUT), .A1 (GND), .A2 (N443));
      NOR2_X1 XNOR_1_3_AND2_NUM251 (.ZN (N1293), .A1 (XNOR_1_1_AND2_NUM251_OUT), .A2 (XNOR_1_2_AND2_NUM251_OUT));
      wire XNOR_1_1_AND2_NUM252_OUT, XNOR_1_2_AND2_NUM252_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM252 (.ZN (XNOR_1_1_AND2_NUM252_OUT), .A1 (N256), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM252 (.ZN (XNOR_1_2_AND2_NUM252_OUT), .A1 (GND), .A2 (N460));
      NOR2_X1 XNOR_1_3_AND2_NUM252 (.ZN (N1296), .A1 (XNOR_1_1_AND2_NUM252_OUT), .A2 (XNOR_1_2_AND2_NUM252_OUT));
      wire XNOR_1_1_AND2_NUM253_OUT, XNOR_1_2_AND2_NUM253_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM253 (.ZN (XNOR_1_1_AND2_NUM253_OUT), .A1 (N256), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM253 (.ZN (XNOR_1_2_AND2_NUM253_OUT), .A1 (GND), .A2 (N477));
      NOR2_X1 XNOR_1_3_AND2_NUM253 (.ZN (N1299), .A1 (XNOR_1_1_AND2_NUM253_OUT), .A2 (XNOR_1_2_AND2_NUM253_OUT));
      wire XNOR_1_1_AND2_NUM254_OUT, XNOR_1_2_AND2_NUM254_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM254 (.ZN (XNOR_1_1_AND2_NUM254_OUT), .A1 (N256), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM254 (.ZN (XNOR_1_2_AND2_NUM254_OUT), .A1 (GND), .A2 (N494));
      NOR2_X1 XNOR_1_3_AND2_NUM254 (.ZN (N1302), .A1 (XNOR_1_1_AND2_NUM254_OUT), .A2 (XNOR_1_2_AND2_NUM254_OUT));
      wire XNOR_1_1_AND2_NUM255_OUT, XNOR_1_2_AND2_NUM255_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM255 (.ZN (XNOR_1_1_AND2_NUM255_OUT), .A1 (N256), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM255 (.ZN (XNOR_1_2_AND2_NUM255_OUT), .A1 (GND), .A2 (N511));
      NOR2_X1 XNOR_1_3_AND2_NUM255 (.ZN (N1305), .A1 (XNOR_1_1_AND2_NUM255_OUT), .A2 (XNOR_1_2_AND2_NUM255_OUT));
      wire XNOR_1_1_AND2_NUM256_OUT, XNOR_1_2_AND2_NUM256_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM256 (.ZN (XNOR_1_1_AND2_NUM256_OUT), .A1 (N256), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM256 (.ZN (XNOR_1_2_AND2_NUM256_OUT), .A1 (GND), .A2 (N528));
      NOR2_X1 XNOR_1_3_AND2_NUM256 (.ZN (N1308), .A1 (XNOR_1_1_AND2_NUM256_OUT), .A2 (XNOR_1_2_AND2_NUM256_OUT));
      NOR2_X1 XNOR_NOT1_NUM257 (.ZN (N1311), .A1 (N591), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM258 (.ZN (N1315), .A1 (N639), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM259 (.ZN (N1319), .A1 (N687), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM260 (.ZN (N1323), .A1 (N735), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM261 (.ZN (N1327), .A1 (N783), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM262 (.ZN (N1331), .A1 (N831), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM263 (.ZN (N1335), .A1 (N879), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM264 (.ZN (N1339), .A1 (N927), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM265 (.ZN (N1343), .A1 (N975), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM266 (.ZN (N1347), .A1 (N1023), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM267 (.ZN (N1351), .A1 (N1071), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM268 (.ZN (N1355), .A1 (N1119), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM269 (.ZN (N1359), .A1 (N1167), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM270 (.ZN (N1363), .A1 (N1215), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM271 (.ZN (N1367), .A1 (N1263), .A2 (GND));
      NOR2_X1 XNOR_NOR2_NUM272 (.ZN (N1371), .A1 (N591), .A2 (N1311));
      NOR2_X1 XNOR_NOT1_NUM273 (.ZN (N1372), .A1 (N1311), .A2 (GND));
      NOR2_X1 XNOR_NOR2_NUM274 (.ZN (N1373), .A1 (N639), .A2 (N1315));
      NOR2_X1 XNOR_NOT1_NUM275 (.ZN (N1374), .A1 (N1315), .A2 (GND));
      NOR2_X1 XNOR_NOR2_NUM276 (.ZN (N1375), .A1 (N687), .A2 (N1319));
      NOR2_X1 XNOR_NOT1_NUM277 (.ZN (N1376), .A1 (N1319), .A2 (GND));
      NOR2_X1 XNOR_NOR2_NUM278 (.ZN (N1377), .A1 (N735), .A2 (N1323));
      NOR2_X1 XNOR_NOT1_NUM279 (.ZN (N1378), .A1 (N1323), .A2 (GND));
      NOR2_X1 XNOR_NOR2_NUM280 (.ZN (N1379), .A1 (N783), .A2 (N1327));
      NOR2_X1 XNOR_NOT1_NUM281 (.ZN (N1380), .A1 (N1327), .A2 (GND));
      NOR2_X1 XNOR_NOR2_NUM282 (.ZN (N1381), .A1 (N831), .A2 (N1331));
      NOR2_X1 XNOR_NOT1_NUM283 (.ZN (N1382), .A1 (N1331), .A2 (GND));
      NOR2_X1 XNOR_NOR2_NUM284 (.ZN (N1383), .A1 (N879), .A2 (N1335));
      NOR2_X1 XNOR_NOT1_NUM285 (.ZN (N1384), .A1 (N1335), .A2 (GND));
      NOR2_X1 XNOR_NOR2_NUM286 (.ZN (N1385), .A1 (N927), .A2 (N1339));
      NOR2_X1 XNOR_NOT1_NUM287 (.ZN (N1386), .A1 (N1339), .A2 (GND));
      NOR2_X1 XNOR_NOR2_NUM288 (.ZN (N1387), .A1 (N975), .A2 (N1343));
      NOR2_X1 XNOR_NOT1_NUM289 (.ZN (N1388), .A1 (N1343), .A2 (GND));
      NOR2_X1 XNOR_NOR2_NUM290 (.ZN (N1389), .A1 (N1023), .A2 (N1347));
      NOR2_X1 XNOR_NOT1_NUM291 (.ZN (N1390), .A1 (N1347), .A2 (GND));
      NOR2_X1 XNOR_NOR2_NUM292 (.ZN (N1391), .A1 (N1071), .A2 (N1351));
      NOR2_X1 XNOR_NOT1_NUM293 (.ZN (N1392), .A1 (N1351), .A2 (GND));
      NOR2_X1 XNOR_NOR2_NUM294 (.ZN (N1393), .A1 (N1119), .A2 (N1355));
      NOR2_X1 XNOR_NOT1_NUM295 (.ZN (N1394), .A1 (N1355), .A2 (GND));
      NOR2_X1 XNOR_NOR2_NUM296 (.ZN (N1395), .A1 (N1167), .A2 (N1359));
      NOR2_X1 XNOR_NOT1_NUM297 (.ZN (N1396), .A1 (N1359), .A2 (GND));
      NOR2_X1 XNOR_NOR2_NUM298 (.ZN (N1397), .A1 (N1215), .A2 (N1363));
      NOR2_X1 XNOR_NOT1_NUM299 (.ZN (N1398), .A1 (N1363), .A2 (GND));
      NOR2_X1 XNOR_NOR2_NUM300 (.ZN (N1399), .A1 (N1263), .A2 (N1367));
      NOR2_X1 XNOR_NOT1_NUM301 (.ZN (N1400), .A1 (N1367), .A2 (GND));
      NOR2_X1 XNOR_NOR2_NUM302 (.ZN (N1401), .A1 (N1371), .A2 (N1372));
      NOR2_X1 XNOR_NOR2_NUM303 (.ZN (N1404), .A1 (N1373), .A2 (N1374));
      NOR2_X1 XNOR_NOR2_NUM304 (.ZN (N1407), .A1 (N1375), .A2 (N1376));
      NOR2_X1 XNOR_NOR2_NUM305 (.ZN (N1410), .A1 (N1377), .A2 (N1378));
      NOR2_X1 XNOR_NOR2_NUM306 (.ZN (N1413), .A1 (N1379), .A2 (N1380));
      NOR2_X1 XNOR_NOR2_NUM307 (.ZN (N1416), .A1 (N1381), .A2 (N1382));
      NOR2_X1 XNOR_NOR2_NUM308 (.ZN (N1419), .A1 (N1383), .A2 (N1384));
      NOR2_X1 XNOR_NOR2_NUM309 (.ZN (N1422), .A1 (N1385), .A2 (N1386));
      NOR2_X1 XNOR_NOR2_NUM310 (.ZN (N1425), .A1 (N1387), .A2 (N1388));
      NOR2_X1 XNOR_NOR2_NUM311 (.ZN (N1428), .A1 (N1389), .A2 (N1390));
      NOR2_X1 XNOR_NOR2_NUM312 (.ZN (N1431), .A1 (N1391), .A2 (N1392));
      NOR2_X1 XNOR_NOR2_NUM313 (.ZN (N1434), .A1 (N1393), .A2 (N1394));
      NOR2_X1 XNOR_NOR2_NUM314 (.ZN (N1437), .A1 (N1395), .A2 (N1396));
      NOR2_X1 XNOR_NOR2_NUM315 (.ZN (N1440), .A1 (N1397), .A2 (N1398));
      NOR2_X1 XNOR_NOR2_NUM316 (.ZN (N1443), .A1 (N1399), .A2 (N1400));
      NOR2_X1 XNOR_NOR2_NUM317 (.ZN (N1446), .A1 (N1401), .A2 (N546));
      NOR2_X1 XNOR_NOR2_NUM318 (.ZN (N1450), .A1 (N1404), .A2 (N594));
      NOR2_X1 XNOR_NOR2_NUM319 (.ZN (N1454), .A1 (N1407), .A2 (N642));
      NOR2_X1 XNOR_NOR2_NUM320 (.ZN (N1458), .A1 (N1410), .A2 (N690));
      NOR2_X1 XNOR_NOR2_NUM321 (.ZN (N1462), .A1 (N1413), .A2 (N738));
      NOR2_X1 XNOR_NOR2_NUM322 (.ZN (N1466), .A1 (N1416), .A2 (N786));
      NOR2_X1 XNOR_NOR2_NUM323 (.ZN (N1470), .A1 (N1419), .A2 (N834));
      NOR2_X1 XNOR_NOR2_NUM324 (.ZN (N1474), .A1 (N1422), .A2 (N882));
      NOR2_X1 XNOR_NOR2_NUM325 (.ZN (N1478), .A1 (N1425), .A2 (N930));
      NOR2_X1 XNOR_NOR2_NUM326 (.ZN (N1482), .A1 (N1428), .A2 (N978));
      NOR2_X1 XNOR_NOR2_NUM327 (.ZN (N1486), .A1 (N1431), .A2 (N1026));
      NOR2_X1 XNOR_NOR2_NUM328 (.ZN (N1490), .A1 (N1434), .A2 (N1074));
      NOR2_X1 XNOR_NOR2_NUM329 (.ZN (N1494), .A1 (N1437), .A2 (N1122));
      NOR2_X1 XNOR_NOR2_NUM330 (.ZN (N1498), .A1 (N1440), .A2 (N1170));
      NOR2_X1 XNOR_NOR2_NUM331 (.ZN (N1502), .A1 (N1443), .A2 (N1218));
      NOR2_X1 XNOR_NOR2_NUM332 (.ZN (N1506), .A1 (N1401), .A2 (N1446));
      NOR2_X1 XNOR_NOR2_NUM333 (.ZN (N1507), .A1 (N1446), .A2 (N546));
      NOR2_X1 XNOR_NOR2_NUM334 (.ZN (N1508), .A1 (N1311), .A2 (N1446));
      NOR2_X1 XNOR_NOR2_NUM335 (.ZN (N1511), .A1 (N1404), .A2 (N1450));
      NOR2_X1 XNOR_NOR2_NUM336 (.ZN (N1512), .A1 (N1450), .A2 (N594));
      NOR2_X1 XNOR_NOR2_NUM337 (.ZN (N1513), .A1 (N1315), .A2 (N1450));
      NOR2_X1 XNOR_NOR2_NUM338 (.ZN (N1516), .A1 (N1407), .A2 (N1454));
      NOR2_X1 XNOR_NOR2_NUM339 (.ZN (N1517), .A1 (N1454), .A2 (N642));
      NOR2_X1 XNOR_NOR2_NUM340 (.ZN (N1518), .A1 (N1319), .A2 (N1454));
      NOR2_X1 XNOR_NOR2_NUM341 (.ZN (N1521), .A1 (N1410), .A2 (N1458));
      NOR2_X1 XNOR_NOR2_NUM342 (.ZN (N1522), .A1 (N1458), .A2 (N690));
      NOR2_X1 XNOR_NOR2_NUM343 (.ZN (N1523), .A1 (N1323), .A2 (N1458));
      NOR2_X1 XNOR_NOR2_NUM344 (.ZN (N1526), .A1 (N1413), .A2 (N1462));
      NOR2_X1 XNOR_NOR2_NUM345 (.ZN (N1527), .A1 (N1462), .A2 (N738));
      NOR2_X1 XNOR_NOR2_NUM346 (.ZN (N1528), .A1 (N1327), .A2 (N1462));
      NOR2_X1 XNOR_NOR2_NUM347 (.ZN (N1531), .A1 (N1416), .A2 (N1466));
      NOR2_X1 XNOR_NOR2_NUM348 (.ZN (N1532), .A1 (N1466), .A2 (N786));
      NOR2_X1 XNOR_NOR2_NUM349 (.ZN (N1533), .A1 (N1331), .A2 (N1466));
      NOR2_X1 XNOR_NOR2_NUM350 (.ZN (N1536), .A1 (N1419), .A2 (N1470));
      NOR2_X1 XNOR_NOR2_NUM351 (.ZN (N1537), .A1 (N1470), .A2 (N834));
      NOR2_X1 XNOR_NOR2_NUM352 (.ZN (N1538), .A1 (N1335), .A2 (N1470));
      NOR2_X1 XNOR_NOR2_NUM353 (.ZN (N1541), .A1 (N1422), .A2 (N1474));
      NOR2_X1 XNOR_NOR2_NUM354 (.ZN (N1542), .A1 (N1474), .A2 (N882));
      NOR2_X1 XNOR_NOR2_NUM355 (.ZN (N1543), .A1 (N1339), .A2 (N1474));
      NOR2_X1 XNOR_NOR2_NUM356 (.ZN (N1546), .A1 (N1425), .A2 (N1478));
      NOR2_X1 XNOR_NOR2_NUM357 (.ZN (N1547), .A1 (N1478), .A2 (N930));
      NOR2_X1 XNOR_NOR2_NUM358 (.ZN (N1548), .A1 (N1343), .A2 (N1478));
      NOR2_X1 XNOR_NOR2_NUM359 (.ZN (N1551), .A1 (N1428), .A2 (N1482));
      NOR2_X1 XNOR_NOR2_NUM360 (.ZN (N1552), .A1 (N1482), .A2 (N978));
      NOR2_X1 XNOR_NOR2_NUM361 (.ZN (N1553), .A1 (N1347), .A2 (N1482));
      NOR2_X1 XNOR_NOR2_NUM362 (.ZN (N1556), .A1 (N1431), .A2 (N1486));
      NOR2_X1 XNOR_NOR2_NUM363 (.ZN (N1557), .A1 (N1486), .A2 (N1026));
      NOR2_X1 XNOR_NOR2_NUM364 (.ZN (N1558), .A1 (N1351), .A2 (N1486));
      NOR2_X1 XNOR_NOR2_NUM365 (.ZN (N1561), .A1 (N1434), .A2 (N1490));
      NOR2_X1 XNOR_NOR2_NUM366 (.ZN (N1562), .A1 (N1490), .A2 (N1074));
      NOR2_X1 XNOR_NOR2_NUM367 (.ZN (N1563), .A1 (N1355), .A2 (N1490));
      NOR2_X1 XNOR_NOR2_NUM368 (.ZN (N1566), .A1 (N1437), .A2 (N1494));
      NOR2_X1 XNOR_NOR2_NUM369 (.ZN (N1567), .A1 (N1494), .A2 (N1122));
      NOR2_X1 XNOR_NOR2_NUM370 (.ZN (N1568), .A1 (N1359), .A2 (N1494));
      NOR2_X1 XNOR_NOR2_NUM371 (.ZN (N1571), .A1 (N1440), .A2 (N1498));
      NOR2_X1 XNOR_NOR2_NUM372 (.ZN (N1572), .A1 (N1498), .A2 (N1170));
      NOR2_X1 XNOR_NOR2_NUM373 (.ZN (N1573), .A1 (N1363), .A2 (N1498));
      NOR2_X1 XNOR_NOR2_NUM374 (.ZN (N1576), .A1 (N1443), .A2 (N1502));
      NOR2_X1 XNOR_NOR2_NUM375 (.ZN (N1577), .A1 (N1502), .A2 (N1218));
      NOR2_X1 XNOR_NOR2_NUM376 (.ZN (N1578), .A1 (N1367), .A2 (N1502));
      NOR2_X1 XNOR_NOR2_NUM377 (.ZN (N1581), .A1 (N1506), .A2 (N1507));
      NOR2_X1 XNOR_NOR2_NUM378 (.ZN (N1582), .A1 (N1511), .A2 (N1512));
      NOR2_X1 XNOR_NOR2_NUM379 (.ZN (N1585), .A1 (N1516), .A2 (N1517));
      NOR2_X1 XNOR_NOR2_NUM380 (.ZN (N1588), .A1 (N1521), .A2 (N1522));
      NOR2_X1 XNOR_NOR2_NUM381 (.ZN (N1591), .A1 (N1526), .A2 (N1527));
      NOR2_X1 XNOR_NOR2_NUM382 (.ZN (N1594), .A1 (N1531), .A2 (N1532));
      NOR2_X1 XNOR_NOR2_NUM383 (.ZN (N1597), .A1 (N1536), .A2 (N1537));
      NOR2_X1 XNOR_NOR2_NUM384 (.ZN (N1600), .A1 (N1541), .A2 (N1542));
      NOR2_X1 XNOR_NOR2_NUM385 (.ZN (N1603), .A1 (N1546), .A2 (N1547));
      NOR2_X1 XNOR_NOR2_NUM386 (.ZN (N1606), .A1 (N1551), .A2 (N1552));
      NOR2_X1 XNOR_NOR2_NUM387 (.ZN (N1609), .A1 (N1556), .A2 (N1557));
      NOR2_X1 XNOR_NOR2_NUM388 (.ZN (N1612), .A1 (N1561), .A2 (N1562));
      NOR2_X1 XNOR_NOR2_NUM389 (.ZN (N1615), .A1 (N1566), .A2 (N1567));
      NOR2_X1 XNOR_NOR2_NUM390 (.ZN (N1618), .A1 (N1571), .A2 (N1572));
      NOR2_X1 XNOR_NOR2_NUM391 (.ZN (N1621), .A1 (N1576), .A2 (N1577));
      NOR2_X1 XNOR_NOR2_NUM392 (.ZN (N1624), .A1 (N1266), .A2 (N1578));
      NOR2_X1 XNOR_NOR2_NUM393 (.ZN (N1628), .A1 (N1582), .A2 (N1508));
      NOR2_X1 XNOR_NOR2_NUM394 (.ZN (N1632), .A1 (N1585), .A2 (N1513));
      NOR2_X1 XNOR_NOR2_NUM395 (.ZN (N1636), .A1 (N1588), .A2 (N1518));
      NOR2_X1 XNOR_NOR2_NUM396 (.ZN (N1640), .A1 (N1591), .A2 (N1523));
      NOR2_X1 XNOR_NOR2_NUM397 (.ZN (N1644), .A1 (N1594), .A2 (N1528));
      NOR2_X1 XNOR_NOR2_NUM398 (.ZN (N1648), .A1 (N1597), .A2 (N1533));
      NOR2_X1 XNOR_NOR2_NUM399 (.ZN (N1652), .A1 (N1600), .A2 (N1538));
      NOR2_X1 XNOR_NOR2_NUM400 (.ZN (N1656), .A1 (N1603), .A2 (N1543));
      NOR2_X1 XNOR_NOR2_NUM401 (.ZN (N1660), .A1 (N1606), .A2 (N1548));
      NOR2_X1 XNOR_NOR2_NUM402 (.ZN (N1664), .A1 (N1609), .A2 (N1553));
      NOR2_X1 XNOR_NOR2_NUM403 (.ZN (N1668), .A1 (N1612), .A2 (N1558));
      NOR2_X1 XNOR_NOR2_NUM404 (.ZN (N1672), .A1 (N1615), .A2 (N1563));
      NOR2_X1 XNOR_NOR2_NUM405 (.ZN (N1676), .A1 (N1618), .A2 (N1568));
      NOR2_X1 XNOR_NOR2_NUM406 (.ZN (N1680), .A1 (N1621), .A2 (N1573));
      NOR2_X1 XNOR_NOR2_NUM407 (.ZN (N1684), .A1 (N1266), .A2 (N1624));
      NOR2_X1 XNOR_NOR2_NUM408 (.ZN (N1685), .A1 (N1624), .A2 (N1578));
      NOR2_X1 XNOR_NOR2_NUM409 (.ZN (N1686), .A1 (N1582), .A2 (N1628));
      NOR2_X1 XNOR_NOR2_NUM410 (.ZN (N1687), .A1 (N1628), .A2 (N1508));
      NOR2_X1 XNOR_NOR2_NUM411 (.ZN (N1688), .A1 (N1585), .A2 (N1632));
      NOR2_X1 XNOR_NOR2_NUM412 (.ZN (N1689), .A1 (N1632), .A2 (N1513));
      NOR2_X1 XNOR_NOR2_NUM413 (.ZN (N1690), .A1 (N1588), .A2 (N1636));
      NOR2_X1 XNOR_NOR2_NUM414 (.ZN (N1691), .A1 (N1636), .A2 (N1518));
      NOR2_X1 XNOR_NOR2_NUM415 (.ZN (N1692), .A1 (N1591), .A2 (N1640));
      NOR2_X1 XNOR_NOR2_NUM416 (.ZN (N1693), .A1 (N1640), .A2 (N1523));
      NOR2_X1 XNOR_NOR2_NUM417 (.ZN (N1694), .A1 (N1594), .A2 (N1644));
      NOR2_X1 XNOR_NOR2_NUM418 (.ZN (N1695), .A1 (N1644), .A2 (N1528));
      NOR2_X1 XNOR_NOR2_NUM419 (.ZN (N1696), .A1 (N1597), .A2 (N1648));
      NOR2_X1 XNOR_NOR2_NUM420 (.ZN (N1697), .A1 (N1648), .A2 (N1533));
      NOR2_X1 XNOR_NOR2_NUM421 (.ZN (N1698), .A1 (N1600), .A2 (N1652));
      NOR2_X1 XNOR_NOR2_NUM422 (.ZN (N1699), .A1 (N1652), .A2 (N1538));
      NOR2_X1 XNOR_NOR2_NUM423 (.ZN (N1700), .A1 (N1603), .A2 (N1656));
      NOR2_X1 XNOR_NOR2_NUM424 (.ZN (N1701), .A1 (N1656), .A2 (N1543));
      NOR2_X1 XNOR_NOR2_NUM425 (.ZN (N1702), .A1 (N1606), .A2 (N1660));
      NOR2_X1 XNOR_NOR2_NUM426 (.ZN (N1703), .A1 (N1660), .A2 (N1548));
      NOR2_X1 XNOR_NOR2_NUM427 (.ZN (N1704), .A1 (N1609), .A2 (N1664));
      NOR2_X1 XNOR_NOR2_NUM428 (.ZN (N1705), .A1 (N1664), .A2 (N1553));
      NOR2_X1 XNOR_NOR2_NUM429 (.ZN (N1706), .A1 (N1612), .A2 (N1668));
      NOR2_X1 XNOR_NOR2_NUM430 (.ZN (N1707), .A1 (N1668), .A2 (N1558));
      NOR2_X1 XNOR_NOR2_NUM431 (.ZN (N1708), .A1 (N1615), .A2 (N1672));
      NOR2_X1 XNOR_NOR2_NUM432 (.ZN (N1709), .A1 (N1672), .A2 (N1563));
      NOR2_X1 XNOR_NOR2_NUM433 (.ZN (N1710), .A1 (N1618), .A2 (N1676));
      NOR2_X1 XNOR_NOR2_NUM434 (.ZN (N1711), .A1 (N1676), .A2 (N1568));
      NOR2_X1 XNOR_NOR2_NUM435 (.ZN (N1712), .A1 (N1621), .A2 (N1680));
      NOR2_X1 XNOR_NOR2_NUM436 (.ZN (N1713), .A1 (N1680), .A2 (N1573));
      NOR2_X1 XNOR_NOR2_NUM437 (.ZN (N1714), .A1 (N1684), .A2 (N1685));
      NOR2_X1 XNOR_NOR2_NUM438 (.ZN (N1717), .A1 (N1686), .A2 (N1687));
      NOR2_X1 XNOR_NOR2_NUM439 (.ZN (N1720), .A1 (N1688), .A2 (N1689));
      NOR2_X1 XNOR_NOR2_NUM440 (.ZN (N1723), .A1 (N1690), .A2 (N1691));
      NOR2_X1 XNOR_NOR2_NUM441 (.ZN (N1726), .A1 (N1692), .A2 (N1693));
      NOR2_X1 XNOR_NOR2_NUM442 (.ZN (N1729), .A1 (N1694), .A2 (N1695));
      NOR2_X1 XNOR_NOR2_NUM443 (.ZN (N1732), .A1 (N1696), .A2 (N1697));
      NOR2_X1 XNOR_NOR2_NUM444 (.ZN (N1735), .A1 (N1698), .A2 (N1699));
      NOR2_X1 XNOR_NOR2_NUM445 (.ZN (N1738), .A1 (N1700), .A2 (N1701));
      NOR2_X1 XNOR_NOR2_NUM446 (.ZN (N1741), .A1 (N1702), .A2 (N1703));
      NOR2_X1 XNOR_NOR2_NUM447 (.ZN (N1744), .A1 (N1704), .A2 (N1705));
      NOR2_X1 XNOR_NOR2_NUM448 (.ZN (N1747), .A1 (N1706), .A2 (N1707));
      NOR2_X1 XNOR_NOR2_NUM449 (.ZN (N1750), .A1 (N1708), .A2 (N1709));
      NOR2_X1 XNOR_NOR2_NUM450 (.ZN (N1753), .A1 (N1710), .A2 (N1711));
      NOR2_X1 XNOR_NOR2_NUM451 (.ZN (N1756), .A1 (N1712), .A2 (N1713));
      NOR2_X1 XNOR_NOR2_NUM452 (.ZN (N1759), .A1 (N1714), .A2 (N1221));
      NOR2_X1 XNOR_NOR2_NUM453 (.ZN (N1763), .A1 (N1717), .A2 (N549));
      NOR2_X1 XNOR_NOR2_NUM454 (.ZN (N1767), .A1 (N1720), .A2 (N597));
      NOR2_X1 XNOR_NOR2_NUM455 (.ZN (N1771), .A1 (N1723), .A2 (N645));
      NOR2_X1 XNOR_NOR2_NUM456 (.ZN (N1775), .A1 (N1726), .A2 (N693));
      NOR2_X1 XNOR_NOR2_NUM457 (.ZN (N1779), .A1 (N1729), .A2 (N741));
      NOR2_X1 XNOR_NOR2_NUM458 (.ZN (N1783), .A1 (N1732), .A2 (N789));
      NOR2_X1 XNOR_NOR2_NUM459 (.ZN (N1787), .A1 (N1735), .A2 (N837));
      NOR2_X1 XNOR_NOR2_NUM460 (.ZN (N1791), .A1 (N1738), .A2 (N885));
      NOR2_X1 XNOR_NOR2_NUM461 (.ZN (N1795), .A1 (N1741), .A2 (N933));
      NOR2_X1 XNOR_NOR2_NUM462 (.ZN (N1799), .A1 (N1744), .A2 (N981));
      NOR2_X1 XNOR_NOR2_NUM463 (.ZN (N1803), .A1 (N1747), .A2 (N1029));
      NOR2_X1 XNOR_NOR2_NUM464 (.ZN (N1807), .A1 (N1750), .A2 (N1077));
      NOR2_X1 XNOR_NOR2_NUM465 (.ZN (N1811), .A1 (N1753), .A2 (N1125));
      NOR2_X1 XNOR_NOR2_NUM466 (.ZN (N1815), .A1 (N1756), .A2 (N1173));
      NOR2_X1 XNOR_NOR2_NUM467 (.ZN (N1819), .A1 (N1714), .A2 (N1759));
      NOR2_X1 XNOR_NOR2_NUM468 (.ZN (N1820), .A1 (N1759), .A2 (N1221));
      NOR2_X1 XNOR_NOR2_NUM469 (.ZN (N1821), .A1 (N1624), .A2 (N1759));
      NOR2_X1 XNOR_NOR2_NUM470 (.ZN (N1824), .A1 (N1717), .A2 (N1763));
      NOR2_X1 XNOR_NOR2_NUM471 (.ZN (N1825), .A1 (N1763), .A2 (N549));
      NOR2_X1 XNOR_NOR2_NUM472 (.ZN (N1826), .A1 (N1628), .A2 (N1763));
      NOR2_X1 XNOR_NOR2_NUM473 (.ZN (N1829), .A1 (N1720), .A2 (N1767));
      NOR2_X1 XNOR_NOR2_NUM474 (.ZN (N1830), .A1 (N1767), .A2 (N597));
      NOR2_X1 XNOR_NOR2_NUM475 (.ZN (N1831), .A1 (N1632), .A2 (N1767));
      NOR2_X1 XNOR_NOR2_NUM476 (.ZN (N1834), .A1 (N1723), .A2 (N1771));
      NOR2_X1 XNOR_NOR2_NUM477 (.ZN (N1835), .A1 (N1771), .A2 (N645));
      NOR2_X1 XNOR_NOR2_NUM478 (.ZN (N1836), .A1 (N1636), .A2 (N1771));
      NOR2_X1 XNOR_NOR2_NUM479 (.ZN (N1839), .A1 (N1726), .A2 (N1775));
      NOR2_X1 XNOR_NOR2_NUM480 (.ZN (N1840), .A1 (N1775), .A2 (N693));
      NOR2_X1 XNOR_NOR2_NUM481 (.ZN (N1841), .A1 (N1640), .A2 (N1775));
      NOR2_X1 XNOR_NOR2_NUM482 (.ZN (N1844), .A1 (N1729), .A2 (N1779));
      NOR2_X1 XNOR_NOR2_NUM483 (.ZN (N1845), .A1 (N1779), .A2 (N741));
      NOR2_X1 XNOR_NOR2_NUM484 (.ZN (N1846), .A1 (N1644), .A2 (N1779));
      NOR2_X1 XNOR_NOR2_NUM485 (.ZN (N1849), .A1 (N1732), .A2 (N1783));
      NOR2_X1 XNOR_NOR2_NUM486 (.ZN (N1850), .A1 (N1783), .A2 (N789));
      NOR2_X1 XNOR_NOR2_NUM487 (.ZN (N1851), .A1 (N1648), .A2 (N1783));
      NOR2_X1 XNOR_NOR2_NUM488 (.ZN (N1854), .A1 (N1735), .A2 (N1787));
      NOR2_X1 XNOR_NOR2_NUM489 (.ZN (N1855), .A1 (N1787), .A2 (N837));
      NOR2_X1 XNOR_NOR2_NUM490 (.ZN (N1856), .A1 (N1652), .A2 (N1787));
      NOR2_X1 XNOR_NOR2_NUM491 (.ZN (N1859), .A1 (N1738), .A2 (N1791));
      NOR2_X1 XNOR_NOR2_NUM492 (.ZN (N1860), .A1 (N1791), .A2 (N885));
      NOR2_X1 XNOR_NOR2_NUM493 (.ZN (N1861), .A1 (N1656), .A2 (N1791));
      NOR2_X1 XNOR_NOR2_NUM494 (.ZN (N1864), .A1 (N1741), .A2 (N1795));
      NOR2_X1 XNOR_NOR2_NUM495 (.ZN (N1865), .A1 (N1795), .A2 (N933));
      NOR2_X1 XNOR_NOR2_NUM496 (.ZN (N1866), .A1 (N1660), .A2 (N1795));
      NOR2_X1 XNOR_NOR2_NUM497 (.ZN (N1869), .A1 (N1744), .A2 (N1799));
      NOR2_X1 XNOR_NOR2_NUM498 (.ZN (N1870), .A1 (N1799), .A2 (N981));
      NOR2_X1 XNOR_NOR2_NUM499 (.ZN (N1871), .A1 (N1664), .A2 (N1799));
      NOR2_X1 XNOR_NOR2_NUM500 (.ZN (N1874), .A1 (N1747), .A2 (N1803));
      NOR2_X1 XNOR_NOR2_NUM501 (.ZN (N1875), .A1 (N1803), .A2 (N1029));
      NOR2_X1 XNOR_NOR2_NUM502 (.ZN (N1876), .A1 (N1668), .A2 (N1803));
      NOR2_X1 XNOR_NOR2_NUM503 (.ZN (N1879), .A1 (N1750), .A2 (N1807));
      NOR2_X1 XNOR_NOR2_NUM504 (.ZN (N1880), .A1 (N1807), .A2 (N1077));
      NOR2_X1 XNOR_NOR2_NUM505 (.ZN (N1881), .A1 (N1672), .A2 (N1807));
      NOR2_X1 XNOR_NOR2_NUM506 (.ZN (N1884), .A1 (N1753), .A2 (N1811));
      NOR2_X1 XNOR_NOR2_NUM507 (.ZN (N1885), .A1 (N1811), .A2 (N1125));
      NOR2_X1 XNOR_NOR2_NUM508 (.ZN (N1886), .A1 (N1676), .A2 (N1811));
      NOR2_X1 XNOR_NOR2_NUM509 (.ZN (N1889), .A1 (N1756), .A2 (N1815));
      NOR2_X1 XNOR_NOR2_NUM510 (.ZN (N1890), .A1 (N1815), .A2 (N1173));
      NOR2_X1 XNOR_NOR2_NUM511 (.ZN (N1891), .A1 (N1680), .A2 (N1815));
      NOR2_X1 XNOR_NOR2_NUM512 (.ZN (N1894), .A1 (N1819), .A2 (N1820));
      NOR2_X1 XNOR_NOR2_NUM513 (.ZN (N1897), .A1 (N1269), .A2 (N1821));
      NOR2_X1 XNOR_NOR2_NUM514 (.ZN (N1901), .A1 (N1824), .A2 (N1825));
      NOR2_X1 XNOR_NOR2_NUM515 (.ZN (N1902), .A1 (N1829), .A2 (N1830));
      NOR2_X1 XNOR_NOR2_NUM516 (.ZN (N1905), .A1 (N1834), .A2 (N1835));
      NOR2_X1 XNOR_NOR2_NUM517 (.ZN (N1908), .A1 (N1839), .A2 (N1840));
      NOR2_X1 XNOR_NOR2_NUM518 (.ZN (N1911), .A1 (N1844), .A2 (N1845));
      NOR2_X1 XNOR_NOR2_NUM519 (.ZN (N1914), .A1 (N1849), .A2 (N1850));
      NOR2_X1 XNOR_NOR2_NUM520 (.ZN (N1917), .A1 (N1854), .A2 (N1855));
      NOR2_X1 XNOR_NOR2_NUM521 (.ZN (N1920), .A1 (N1859), .A2 (N1860));
      NOR2_X1 XNOR_NOR2_NUM522 (.ZN (N1923), .A1 (N1864), .A2 (N1865));
      NOR2_X1 XNOR_NOR2_NUM523 (.ZN (N1926), .A1 (N1869), .A2 (N1870));
      NOR2_X1 XNOR_NOR2_NUM524 (.ZN (N1929), .A1 (N1874), .A2 (N1875));
      NOR2_X1 XNOR_NOR2_NUM525 (.ZN (N1932), .A1 (N1879), .A2 (N1880));
      NOR2_X1 XNOR_NOR2_NUM526 (.ZN (N1935), .A1 (N1884), .A2 (N1885));
      NOR2_X1 XNOR_NOR2_NUM527 (.ZN (N1938), .A1 (N1889), .A2 (N1890));
      NOR2_X1 XNOR_NOR2_NUM528 (.ZN (N1941), .A1 (N1894), .A2 (N1891));
      NOR2_X1 XNOR_NOR2_NUM529 (.ZN (N1945), .A1 (N1269), .A2 (N1897));
      NOR2_X1 XNOR_NOR2_NUM530 (.ZN (N1946), .A1 (N1897), .A2 (N1821));
      NOR2_X1 XNOR_NOR2_NUM531 (.ZN (N1947), .A1 (N1902), .A2 (N1826));
      NOR2_X1 XNOR_NOR2_NUM532 (.ZN (N1951), .A1 (N1905), .A2 (N1831));
      NOR2_X1 XNOR_NOR2_NUM533 (.ZN (N1955), .A1 (N1908), .A2 (N1836));
      NOR2_X1 XNOR_NOR2_NUM534 (.ZN (N1959), .A1 (N1911), .A2 (N1841));
      NOR2_X1 XNOR_NOR2_NUM535 (.ZN (N1963), .A1 (N1914), .A2 (N1846));
      NOR2_X1 XNOR_NOR2_NUM536 (.ZN (N1967), .A1 (N1917), .A2 (N1851));
      NOR2_X1 XNOR_NOR2_NUM537 (.ZN (N1971), .A1 (N1920), .A2 (N1856));
      NOR2_X1 XNOR_NOR2_NUM538 (.ZN (N1975), .A1 (N1923), .A2 (N1861));
      NOR2_X1 XNOR_NOR2_NUM539 (.ZN (N1979), .A1 (N1926), .A2 (N1866));
      NOR2_X1 XNOR_NOR2_NUM540 (.ZN (N1983), .A1 (N1929), .A2 (N1871));
      NOR2_X1 XNOR_NOR2_NUM541 (.ZN (N1987), .A1 (N1932), .A2 (N1876));
      NOR2_X1 XNOR_NOR2_NUM542 (.ZN (N1991), .A1 (N1935), .A2 (N1881));
      NOR2_X1 XNOR_NOR2_NUM543 (.ZN (N1995), .A1 (N1938), .A2 (N1886));
      NOR2_X1 XNOR_NOR2_NUM544 (.ZN (N1999), .A1 (N1894), .A2 (N1941));
      NOR2_X1 XNOR_NOR2_NUM545 (.ZN (N2000), .A1 (N1941), .A2 (N1891));
      NOR2_X1 XNOR_NOR2_NUM546 (.ZN (N2001), .A1 (N1945), .A2 (N1946));
      NOR2_X1 XNOR_NOR2_NUM547 (.ZN (N2004), .A1 (N1902), .A2 (N1947));
      NOR2_X1 XNOR_NOR2_NUM548 (.ZN (N2005), .A1 (N1947), .A2 (N1826));
      NOR2_X1 XNOR_NOR2_NUM549 (.ZN (N2006), .A1 (N1905), .A2 (N1951));
      NOR2_X1 XNOR_NOR2_NUM550 (.ZN (N2007), .A1 (N1951), .A2 (N1831));
      NOR2_X1 XNOR_NOR2_NUM551 (.ZN (N2008), .A1 (N1908), .A2 (N1955));
      NOR2_X1 XNOR_NOR2_NUM552 (.ZN (N2009), .A1 (N1955), .A2 (N1836));
      NOR2_X1 XNOR_NOR2_NUM553 (.ZN (N2010), .A1 (N1911), .A2 (N1959));
      NOR2_X1 XNOR_NOR2_NUM554 (.ZN (N2011), .A1 (N1959), .A2 (N1841));
      NOR2_X1 XNOR_NOR2_NUM555 (.ZN (N2012), .A1 (N1914), .A2 (N1963));
      NOR2_X1 XNOR_NOR2_NUM556 (.ZN (N2013), .A1 (N1963), .A2 (N1846));
      NOR2_X1 XNOR_NOR2_NUM557 (.ZN (N2014), .A1 (N1917), .A2 (N1967));
      NOR2_X1 XNOR_NOR2_NUM558 (.ZN (N2015), .A1 (N1967), .A2 (N1851));
      NOR2_X1 XNOR_NOR2_NUM559 (.ZN (N2016), .A1 (N1920), .A2 (N1971));
      NOR2_X1 XNOR_NOR2_NUM560 (.ZN (N2017), .A1 (N1971), .A2 (N1856));
      NOR2_X1 XNOR_NOR2_NUM561 (.ZN (N2018), .A1 (N1923), .A2 (N1975));
      NOR2_X1 XNOR_NOR2_NUM562 (.ZN (N2019), .A1 (N1975), .A2 (N1861));
      NOR2_X1 XNOR_NOR2_NUM563 (.ZN (N2020), .A1 (N1926), .A2 (N1979));
      NOR2_X1 XNOR_NOR2_NUM564 (.ZN (N2021), .A1 (N1979), .A2 (N1866));
      NOR2_X1 XNOR_NOR2_NUM565 (.ZN (N2022), .A1 (N1929), .A2 (N1983));
      NOR2_X1 XNOR_NOR2_NUM566 (.ZN (N2023), .A1 (N1983), .A2 (N1871));
      NOR2_X1 XNOR_NOR2_NUM567 (.ZN (N2024), .A1 (N1932), .A2 (N1987));
      NOR2_X1 XNOR_NOR2_NUM568 (.ZN (N2025), .A1 (N1987), .A2 (N1876));
      NOR2_X1 XNOR_NOR2_NUM569 (.ZN (N2026), .A1 (N1935), .A2 (N1991));
      NOR2_X1 XNOR_NOR2_NUM570 (.ZN (N2027), .A1 (N1991), .A2 (N1881));
      NOR2_X1 XNOR_NOR2_NUM571 (.ZN (N2028), .A1 (N1938), .A2 (N1995));
      NOR2_X1 XNOR_NOR2_NUM572 (.ZN (N2029), .A1 (N1995), .A2 (N1886));
      NOR2_X1 XNOR_NOR2_NUM573 (.ZN (N2030), .A1 (N1999), .A2 (N2000));
      NOR2_X1 XNOR_NOR2_NUM574 (.ZN (N2033), .A1 (N2001), .A2 (N1224));
      NOR2_X1 XNOR_NOR2_NUM575 (.ZN (N2037), .A1 (N2004), .A2 (N2005));
      NOR2_X1 XNOR_NOR2_NUM576 (.ZN (N2040), .A1 (N2006), .A2 (N2007));
      NOR2_X1 XNOR_NOR2_NUM577 (.ZN (N2043), .A1 (N2008), .A2 (N2009));
      NOR2_X1 XNOR_NOR2_NUM578 (.ZN (N2046), .A1 (N2010), .A2 (N2011));
      NOR2_X1 XNOR_NOR2_NUM579 (.ZN (N2049), .A1 (N2012), .A2 (N2013));
      NOR2_X1 XNOR_NOR2_NUM580 (.ZN (N2052), .A1 (N2014), .A2 (N2015));
      NOR2_X1 XNOR_NOR2_NUM581 (.ZN (N2055), .A1 (N2016), .A2 (N2017));
      NOR2_X1 XNOR_NOR2_NUM582 (.ZN (N2058), .A1 (N2018), .A2 (N2019));
      NOR2_X1 XNOR_NOR2_NUM583 (.ZN (N2061), .A1 (N2020), .A2 (N2021));
      NOR2_X1 XNOR_NOR2_NUM584 (.ZN (N2064), .A1 (N2022), .A2 (N2023));
      NOR2_X1 XNOR_NOR2_NUM585 (.ZN (N2067), .A1 (N2024), .A2 (N2025));
      NOR2_X1 XNOR_NOR2_NUM586 (.ZN (N2070), .A1 (N2026), .A2 (N2027));
      NOR2_X1 XNOR_NOR2_NUM587 (.ZN (N2073), .A1 (N2028), .A2 (N2029));
      NOR2_X1 XNOR_NOR2_NUM588 (.ZN (N2076), .A1 (N2030), .A2 (N1176));
      NOR2_X1 XNOR_NOR2_NUM589 (.ZN (N2080), .A1 (N2001), .A2 (N2033));
      NOR2_X1 XNOR_NOR2_NUM590 (.ZN (N2081), .A1 (N2033), .A2 (N1224));
      NOR2_X1 XNOR_NOR2_NUM591 (.ZN (N2082), .A1 (N1897), .A2 (N2033));
      NOR2_X1 XNOR_NOR2_NUM592 (.ZN (N2085), .A1 (N2037), .A2 (N552));
      NOR2_X1 XNOR_NOR2_NUM593 (.ZN (N2089), .A1 (N2040), .A2 (N600));
      NOR2_X1 XNOR_NOR2_NUM594 (.ZN (N2093), .A1 (N2043), .A2 (N648));
      NOR2_X1 XNOR_NOR2_NUM595 (.ZN (N2097), .A1 (N2046), .A2 (N696));
      NOR2_X1 XNOR_NOR2_NUM596 (.ZN (N2101), .A1 (N2049), .A2 (N744));
      NOR2_X1 XNOR_NOR2_NUM597 (.ZN (N2105), .A1 (N2052), .A2 (N792));
      NOR2_X1 XNOR_NOR2_NUM598 (.ZN (N2109), .A1 (N2055), .A2 (N840));
      NOR2_X1 XNOR_NOR2_NUM599 (.ZN (N2113), .A1 (N2058), .A2 (N888));
      NOR2_X1 XNOR_NOR2_NUM600 (.ZN (N2117), .A1 (N2061), .A2 (N936));
      NOR2_X1 XNOR_NOR2_NUM601 (.ZN (N2121), .A1 (N2064), .A2 (N984));
      NOR2_X1 XNOR_NOR2_NUM602 (.ZN (N2125), .A1 (N2067), .A2 (N1032));
      NOR2_X1 XNOR_NOR2_NUM603 (.ZN (N2129), .A1 (N2070), .A2 (N1080));
      NOR2_X1 XNOR_NOR2_NUM604 (.ZN (N2133), .A1 (N2073), .A2 (N1128));
      NOR2_X1 XNOR_NOR2_NUM605 (.ZN (N2137), .A1 (N2030), .A2 (N2076));
      NOR2_X1 XNOR_NOR2_NUM606 (.ZN (N2138), .A1 (N2076), .A2 (N1176));
      NOR2_X1 XNOR_NOR2_NUM607 (.ZN (N2139), .A1 (N1941), .A2 (N2076));
      NOR2_X1 XNOR_NOR2_NUM608 (.ZN (N2142), .A1 (N2080), .A2 (N2081));
      NOR2_X1 XNOR_NOR2_NUM609 (.ZN (N2145), .A1 (N1272), .A2 (N2082));
      NOR2_X1 XNOR_NOR2_NUM610 (.ZN (N2149), .A1 (N2037), .A2 (N2085));
      NOR2_X1 XNOR_NOR2_NUM611 (.ZN (N2150), .A1 (N2085), .A2 (N552));
      NOR2_X1 XNOR_NOR2_NUM612 (.ZN (N2151), .A1 (N1947), .A2 (N2085));
      NOR2_X1 XNOR_NOR2_NUM613 (.ZN (N2154), .A1 (N2040), .A2 (N2089));
      NOR2_X1 XNOR_NOR2_NUM614 (.ZN (N2155), .A1 (N2089), .A2 (N600));
      NOR2_X1 XNOR_NOR2_NUM615 (.ZN (N2156), .A1 (N1951), .A2 (N2089));
      NOR2_X1 XNOR_NOR2_NUM616 (.ZN (N2159), .A1 (N2043), .A2 (N2093));
      NOR2_X1 XNOR_NOR2_NUM617 (.ZN (N2160), .A1 (N2093), .A2 (N648));
      NOR2_X1 XNOR_NOR2_NUM618 (.ZN (N2161), .A1 (N1955), .A2 (N2093));
      NOR2_X1 XNOR_NOR2_NUM619 (.ZN (N2164), .A1 (N2046), .A2 (N2097));
      NOR2_X1 XNOR_NOR2_NUM620 (.ZN (N2165), .A1 (N2097), .A2 (N696));
      NOR2_X1 XNOR_NOR2_NUM621 (.ZN (N2166), .A1 (N1959), .A2 (N2097));
      NOR2_X1 XNOR_NOR2_NUM622 (.ZN (N2169), .A1 (N2049), .A2 (N2101));
      NOR2_X1 XNOR_NOR2_NUM623 (.ZN (N2170), .A1 (N2101), .A2 (N744));
      NOR2_X1 XNOR_NOR2_NUM624 (.ZN (N2171), .A1 (N1963), .A2 (N2101));
      NOR2_X1 XNOR_NOR2_NUM625 (.ZN (N2174), .A1 (N2052), .A2 (N2105));
      NOR2_X1 XNOR_NOR2_NUM626 (.ZN (N2175), .A1 (N2105), .A2 (N792));
      NOR2_X1 XNOR_NOR2_NUM627 (.ZN (N2176), .A1 (N1967), .A2 (N2105));
      NOR2_X1 XNOR_NOR2_NUM628 (.ZN (N2179), .A1 (N2055), .A2 (N2109));
      NOR2_X1 XNOR_NOR2_NUM629 (.ZN (N2180), .A1 (N2109), .A2 (N840));
      NOR2_X1 XNOR_NOR2_NUM630 (.ZN (N2181), .A1 (N1971), .A2 (N2109));
      NOR2_X1 XNOR_NOR2_NUM631 (.ZN (N2184), .A1 (N2058), .A2 (N2113));
      NOR2_X1 XNOR_NOR2_NUM632 (.ZN (N2185), .A1 (N2113), .A2 (N888));
      NOR2_X1 XNOR_NOR2_NUM633 (.ZN (N2186), .A1 (N1975), .A2 (N2113));
      NOR2_X1 XNOR_NOR2_NUM634 (.ZN (N2189), .A1 (N2061), .A2 (N2117));
      NOR2_X1 XNOR_NOR2_NUM635 (.ZN (N2190), .A1 (N2117), .A2 (N936));
      NOR2_X1 XNOR_NOR2_NUM636 (.ZN (N2191), .A1 (N1979), .A2 (N2117));
      NOR2_X1 XNOR_NOR2_NUM637 (.ZN (N2194), .A1 (N2064), .A2 (N2121));
      NOR2_X1 XNOR_NOR2_NUM638 (.ZN (N2195), .A1 (N2121), .A2 (N984));
      NOR2_X1 XNOR_NOR2_NUM639 (.ZN (N2196), .A1 (N1983), .A2 (N2121));
      NOR2_X1 XNOR_NOR2_NUM640 (.ZN (N2199), .A1 (N2067), .A2 (N2125));
      NOR2_X1 XNOR_NOR2_NUM641 (.ZN (N2200), .A1 (N2125), .A2 (N1032));
      NOR2_X1 XNOR_NOR2_NUM642 (.ZN (N2201), .A1 (N1987), .A2 (N2125));
      NOR2_X1 XNOR_NOR2_NUM643 (.ZN (N2204), .A1 (N2070), .A2 (N2129));
      NOR2_X1 XNOR_NOR2_NUM644 (.ZN (N2205), .A1 (N2129), .A2 (N1080));
      NOR2_X1 XNOR_NOR2_NUM645 (.ZN (N2206), .A1 (N1991), .A2 (N2129));
      NOR2_X1 XNOR_NOR2_NUM646 (.ZN (N2209), .A1 (N2073), .A2 (N2133));
      NOR2_X1 XNOR_NOR2_NUM647 (.ZN (N2210), .A1 (N2133), .A2 (N1128));
      NOR2_X1 XNOR_NOR2_NUM648 (.ZN (N2211), .A1 (N1995), .A2 (N2133));
      NOR2_X1 XNOR_NOR2_NUM649 (.ZN (N2214), .A1 (N2137), .A2 (N2138));
      NOR2_X1 XNOR_NOR2_NUM650 (.ZN (N2217), .A1 (N2142), .A2 (N2139));
      NOR2_X1 XNOR_NOR2_NUM651 (.ZN (N2221), .A1 (N1272), .A2 (N2145));
      NOR2_X1 XNOR_NOR2_NUM652 (.ZN (N2222), .A1 (N2145), .A2 (N2082));
      NOR2_X1 XNOR_NOR2_NUM653 (.ZN (N2223), .A1 (N2149), .A2 (N2150));
      NOR2_X1 XNOR_NOR2_NUM654 (.ZN (N2224), .A1 (N2154), .A2 (N2155));
      NOR2_X1 XNOR_NOR2_NUM655 (.ZN (N2227), .A1 (N2159), .A2 (N2160));
      NOR2_X1 XNOR_NOR2_NUM656 (.ZN (N2230), .A1 (N2164), .A2 (N2165));
      NOR2_X1 XNOR_NOR2_NUM657 (.ZN (N2233), .A1 (N2169), .A2 (N2170));
      NOR2_X1 XNOR_NOR2_NUM658 (.ZN (N2236), .A1 (N2174), .A2 (N2175));
      NOR2_X1 XNOR_NOR2_NUM659 (.ZN (N2239), .A1 (N2179), .A2 (N2180));
      NOR2_X1 XNOR_NOR2_NUM660 (.ZN (N2242), .A1 (N2184), .A2 (N2185));
      NOR2_X1 XNOR_NOR2_NUM661 (.ZN (N2245), .A1 (N2189), .A2 (N2190));
      NOR2_X1 XNOR_NOR2_NUM662 (.ZN (N2248), .A1 (N2194), .A2 (N2195));
      NOR2_X1 XNOR_NOR2_NUM663 (.ZN (N2251), .A1 (N2199), .A2 (N2200));
      NOR2_X1 XNOR_NOR2_NUM664 (.ZN (N2254), .A1 (N2204), .A2 (N2205));
      NOR2_X1 XNOR_NOR2_NUM665 (.ZN (N2257), .A1 (N2209), .A2 (N2210));
      NOR2_X1 XNOR_NOR2_NUM666 (.ZN (N2260), .A1 (N2214), .A2 (N2211));
      NOR2_X1 XNOR_NOR2_NUM667 (.ZN (N2264), .A1 (N2142), .A2 (N2217));
      NOR2_X1 XNOR_NOR2_NUM668 (.ZN (N2265), .A1 (N2217), .A2 (N2139));
      NOR2_X1 XNOR_NOR2_NUM669 (.ZN (N2266), .A1 (N2221), .A2 (N2222));
      NOR2_X1 XNOR_NOR2_NUM670 (.ZN (N2269), .A1 (N2224), .A2 (N2151));
      NOR2_X1 XNOR_NOR2_NUM671 (.ZN (N2273), .A1 (N2227), .A2 (N2156));
      NOR2_X1 XNOR_NOR2_NUM672 (.ZN (N2277), .A1 (N2230), .A2 (N2161));
      NOR2_X1 XNOR_NOR2_NUM673 (.ZN (N2281), .A1 (N2233), .A2 (N2166));
      NOR2_X1 XNOR_NOR2_NUM674 (.ZN (N2285), .A1 (N2236), .A2 (N2171));
      NOR2_X1 XNOR_NOR2_NUM675 (.ZN (N2289), .A1 (N2239), .A2 (N2176));
      NOR2_X1 XNOR_NOR2_NUM676 (.ZN (N2293), .A1 (N2242), .A2 (N2181));
      NOR2_X1 XNOR_NOR2_NUM677 (.ZN (N2297), .A1 (N2245), .A2 (N2186));
      NOR2_X1 XNOR_NOR2_NUM678 (.ZN (N2301), .A1 (N2248), .A2 (N2191));
      NOR2_X1 XNOR_NOR2_NUM679 (.ZN (N2305), .A1 (N2251), .A2 (N2196));
      NOR2_X1 XNOR_NOR2_NUM680 (.ZN (N2309), .A1 (N2254), .A2 (N2201));
      NOR2_X1 XNOR_NOR2_NUM681 (.ZN (N2313), .A1 (N2257), .A2 (N2206));
      NOR2_X1 XNOR_NOR2_NUM682 (.ZN (N2317), .A1 (N2214), .A2 (N2260));
      NOR2_X1 XNOR_NOR2_NUM683 (.ZN (N2318), .A1 (N2260), .A2 (N2211));
      NOR2_X1 XNOR_NOR2_NUM684 (.ZN (N2319), .A1 (N2264), .A2 (N2265));
      NOR2_X1 XNOR_NOR2_NUM685 (.ZN (N2322), .A1 (N2266), .A2 (N1227));
      NOR2_X1 XNOR_NOR2_NUM686 (.ZN (N2326), .A1 (N2224), .A2 (N2269));
      NOR2_X1 XNOR_NOR2_NUM687 (.ZN (N2327), .A1 (N2269), .A2 (N2151));
      NOR2_X1 XNOR_NOR2_NUM688 (.ZN (N2328), .A1 (N2227), .A2 (N2273));
      NOR2_X1 XNOR_NOR2_NUM689 (.ZN (N2329), .A1 (N2273), .A2 (N2156));
      NOR2_X1 XNOR_NOR2_NUM690 (.ZN (N2330), .A1 (N2230), .A2 (N2277));
      NOR2_X1 XNOR_NOR2_NUM691 (.ZN (N2331), .A1 (N2277), .A2 (N2161));
      NOR2_X1 XNOR_NOR2_NUM692 (.ZN (N2332), .A1 (N2233), .A2 (N2281));
      NOR2_X1 XNOR_NOR2_NUM693 (.ZN (N2333), .A1 (N2281), .A2 (N2166));
      NOR2_X1 XNOR_NOR2_NUM694 (.ZN (N2334), .A1 (N2236), .A2 (N2285));
      NOR2_X1 XNOR_NOR2_NUM695 (.ZN (N2335), .A1 (N2285), .A2 (N2171));
      NOR2_X1 XNOR_NOR2_NUM696 (.ZN (N2336), .A1 (N2239), .A2 (N2289));
      NOR2_X1 XNOR_NOR2_NUM697 (.ZN (N2337), .A1 (N2289), .A2 (N2176));
      NOR2_X1 XNOR_NOR2_NUM698 (.ZN (N2338), .A1 (N2242), .A2 (N2293));
      NOR2_X1 XNOR_NOR2_NUM699 (.ZN (N2339), .A1 (N2293), .A2 (N2181));
      NOR2_X1 XNOR_NOR2_NUM700 (.ZN (N2340), .A1 (N2245), .A2 (N2297));
      NOR2_X1 XNOR_NOR2_NUM701 (.ZN (N2341), .A1 (N2297), .A2 (N2186));
      NOR2_X1 XNOR_NOR2_NUM702 (.ZN (N2342), .A1 (N2248), .A2 (N2301));
      NOR2_X1 XNOR_NOR2_NUM703 (.ZN (N2343), .A1 (N2301), .A2 (N2191));
      NOR2_X1 XNOR_NOR2_NUM704 (.ZN (N2344), .A1 (N2251), .A2 (N2305));
      NOR2_X1 XNOR_NOR2_NUM705 (.ZN (N2345), .A1 (N2305), .A2 (N2196));
      NOR2_X1 XNOR_NOR2_NUM706 (.ZN (N2346), .A1 (N2254), .A2 (N2309));
      NOR2_X1 XNOR_NOR2_NUM707 (.ZN (N2347), .A1 (N2309), .A2 (N2201));
      NOR2_X1 XNOR_NOR2_NUM708 (.ZN (N2348), .A1 (N2257), .A2 (N2313));
      NOR2_X1 XNOR_NOR2_NUM709 (.ZN (N2349), .A1 (N2313), .A2 (N2206));
      NOR2_X1 XNOR_NOR2_NUM710 (.ZN (N2350), .A1 (N2317), .A2 (N2318));
      NOR2_X1 XNOR_NOR2_NUM711 (.ZN (N2353), .A1 (N2319), .A2 (N1179));
      NOR2_X1 XNOR_NOR2_NUM712 (.ZN (N2357), .A1 (N2266), .A2 (N2322));
      NOR2_X1 XNOR_NOR2_NUM713 (.ZN (N2358), .A1 (N2322), .A2 (N1227));
      NOR2_X1 XNOR_NOR2_NUM714 (.ZN (N2359), .A1 (N2145), .A2 (N2322));
      NOR2_X1 XNOR_NOR2_NUM715 (.ZN (N2362), .A1 (N2326), .A2 (N2327));
      NOR2_X1 XNOR_NOR2_NUM716 (.ZN (N2365), .A1 (N2328), .A2 (N2329));
      NOR2_X1 XNOR_NOR2_NUM717 (.ZN (N2368), .A1 (N2330), .A2 (N2331));
      NOR2_X1 XNOR_NOR2_NUM718 (.ZN (N2371), .A1 (N2332), .A2 (N2333));
      NOR2_X1 XNOR_NOR2_NUM719 (.ZN (N2374), .A1 (N2334), .A2 (N2335));
      NOR2_X1 XNOR_NOR2_NUM720 (.ZN (N2377), .A1 (N2336), .A2 (N2337));
      NOR2_X1 XNOR_NOR2_NUM721 (.ZN (N2380), .A1 (N2338), .A2 (N2339));
      NOR2_X1 XNOR_NOR2_NUM722 (.ZN (N2383), .A1 (N2340), .A2 (N2341));
      NOR2_X1 XNOR_NOR2_NUM723 (.ZN (N2386), .A1 (N2342), .A2 (N2343));
      NOR2_X1 XNOR_NOR2_NUM724 (.ZN (N2389), .A1 (N2344), .A2 (N2345));
      NOR2_X1 XNOR_NOR2_NUM725 (.ZN (N2392), .A1 (N2346), .A2 (N2347));
      NOR2_X1 XNOR_NOR2_NUM726 (.ZN (N2395), .A1 (N2348), .A2 (N2349));
      NOR2_X1 XNOR_NOR2_NUM727 (.ZN (N2398), .A1 (N2350), .A2 (N1131));
      NOR2_X1 XNOR_NOR2_NUM728 (.ZN (N2402), .A1 (N2319), .A2 (N2353));
      NOR2_X1 XNOR_NOR2_NUM729 (.ZN (N2403), .A1 (N2353), .A2 (N1179));
      NOR2_X1 XNOR_NOR2_NUM730 (.ZN (N2404), .A1 (N2217), .A2 (N2353));
      NOR2_X1 XNOR_NOR2_NUM731 (.ZN (N2407), .A1 (N2357), .A2 (N2358));
      NOR2_X1 XNOR_NOR2_NUM732 (.ZN (N2410), .A1 (N1275), .A2 (N2359));
      NOR2_X1 XNOR_NOR2_NUM733 (.ZN (N2414), .A1 (N2362), .A2 (N555));
      NOR2_X1 XNOR_NOR2_NUM734 (.ZN (N2418), .A1 (N2365), .A2 (N603));
      NOR2_X1 XNOR_NOR2_NUM735 (.ZN (N2422), .A1 (N2368), .A2 (N651));
      NOR2_X1 XNOR_NOR2_NUM736 (.ZN (N2426), .A1 (N2371), .A2 (N699));
      NOR2_X1 XNOR_NOR2_NUM737 (.ZN (N2430), .A1 (N2374), .A2 (N747));
      NOR2_X1 XNOR_NOR2_NUM738 (.ZN (N2434), .A1 (N2377), .A2 (N795));
      NOR2_X1 XNOR_NOR2_NUM739 (.ZN (N2438), .A1 (N2380), .A2 (N843));
      NOR2_X1 XNOR_NOR2_NUM740 (.ZN (N2442), .A1 (N2383), .A2 (N891));
      NOR2_X1 XNOR_NOR2_NUM741 (.ZN (N2446), .A1 (N2386), .A2 (N939));
      NOR2_X1 XNOR_NOR2_NUM742 (.ZN (N2450), .A1 (N2389), .A2 (N987));
      NOR2_X1 XNOR_NOR2_NUM743 (.ZN (N2454), .A1 (N2392), .A2 (N1035));
      NOR2_X1 XNOR_NOR2_NUM744 (.ZN (N2458), .A1 (N2395), .A2 (N1083));
      NOR2_X1 XNOR_NOR2_NUM745 (.ZN (N2462), .A1 (N2350), .A2 (N2398));
      NOR2_X1 XNOR_NOR2_NUM746 (.ZN (N2463), .A1 (N2398), .A2 (N1131));
      NOR2_X1 XNOR_NOR2_NUM747 (.ZN (N2464), .A1 (N2260), .A2 (N2398));
      NOR2_X1 XNOR_NOR2_NUM748 (.ZN (N2467), .A1 (N2402), .A2 (N2403));
      NOR2_X1 XNOR_NOR2_NUM749 (.ZN (N2470), .A1 (N2407), .A2 (N2404));
      NOR2_X1 XNOR_NOR2_NUM750 (.ZN (N2474), .A1 (N1275), .A2 (N2410));
      NOR2_X1 XNOR_NOR2_NUM751 (.ZN (N2475), .A1 (N2410), .A2 (N2359));
      NOR2_X1 XNOR_NOR2_NUM752 (.ZN (N2476), .A1 (N2362), .A2 (N2414));
      NOR2_X1 XNOR_NOR2_NUM753 (.ZN (N2477), .A1 (N2414), .A2 (N555));
      NOR2_X1 XNOR_NOR2_NUM754 (.ZN (N2478), .A1 (N2269), .A2 (N2414));
      NOR2_X1 XNOR_NOR2_NUM755 (.ZN (N2481), .A1 (N2365), .A2 (N2418));
      NOR2_X1 XNOR_NOR2_NUM756 (.ZN (N2482), .A1 (N2418), .A2 (N603));
      NOR2_X1 XNOR_NOR2_NUM757 (.ZN (N2483), .A1 (N2273), .A2 (N2418));
      NOR2_X1 XNOR_NOR2_NUM758 (.ZN (N2486), .A1 (N2368), .A2 (N2422));
      NOR2_X1 XNOR_NOR2_NUM759 (.ZN (N2487), .A1 (N2422), .A2 (N651));
      NOR2_X1 XNOR_NOR2_NUM760 (.ZN (N2488), .A1 (N2277), .A2 (N2422));
      NOR2_X1 XNOR_NOR2_NUM761 (.ZN (N2491), .A1 (N2371), .A2 (N2426));
      NOR2_X1 XNOR_NOR2_NUM762 (.ZN (N2492), .A1 (N2426), .A2 (N699));
      NOR2_X1 XNOR_NOR2_NUM763 (.ZN (N2493), .A1 (N2281), .A2 (N2426));
      NOR2_X1 XNOR_NOR2_NUM764 (.ZN (N2496), .A1 (N2374), .A2 (N2430));
      NOR2_X1 XNOR_NOR2_NUM765 (.ZN (N2497), .A1 (N2430), .A2 (N747));
      NOR2_X1 XNOR_NOR2_NUM766 (.ZN (N2498), .A1 (N2285), .A2 (N2430));
      NOR2_X1 XNOR_NOR2_NUM767 (.ZN (N2501), .A1 (N2377), .A2 (N2434));
      NOR2_X1 XNOR_NOR2_NUM768 (.ZN (N2502), .A1 (N2434), .A2 (N795));
      NOR2_X1 XNOR_NOR2_NUM769 (.ZN (N2503), .A1 (N2289), .A2 (N2434));
      NOR2_X1 XNOR_NOR2_NUM770 (.ZN (N2506), .A1 (N2380), .A2 (N2438));
      NOR2_X1 XNOR_NOR2_NUM771 (.ZN (N2507), .A1 (N2438), .A2 (N843));
      NOR2_X1 XNOR_NOR2_NUM772 (.ZN (N2508), .A1 (N2293), .A2 (N2438));
      NOR2_X1 XNOR_NOR2_NUM773 (.ZN (N2511), .A1 (N2383), .A2 (N2442));
      NOR2_X1 XNOR_NOR2_NUM774 (.ZN (N2512), .A1 (N2442), .A2 (N891));
      NOR2_X1 XNOR_NOR2_NUM775 (.ZN (N2513), .A1 (N2297), .A2 (N2442));
      NOR2_X1 XNOR_NOR2_NUM776 (.ZN (N2516), .A1 (N2386), .A2 (N2446));
      NOR2_X1 XNOR_NOR2_NUM777 (.ZN (N2517), .A1 (N2446), .A2 (N939));
      NOR2_X1 XNOR_NOR2_NUM778 (.ZN (N2518), .A1 (N2301), .A2 (N2446));
      NOR2_X1 XNOR_NOR2_NUM779 (.ZN (N2521), .A1 (N2389), .A2 (N2450));
      NOR2_X1 XNOR_NOR2_NUM780 (.ZN (N2522), .A1 (N2450), .A2 (N987));
      NOR2_X1 XNOR_NOR2_NUM781 (.ZN (N2523), .A1 (N2305), .A2 (N2450));
      NOR2_X1 XNOR_NOR2_NUM782 (.ZN (N2526), .A1 (N2392), .A2 (N2454));
      NOR2_X1 XNOR_NOR2_NUM783 (.ZN (N2527), .A1 (N2454), .A2 (N1035));
      NOR2_X1 XNOR_NOR2_NUM784 (.ZN (N2528), .A1 (N2309), .A2 (N2454));
      NOR2_X1 XNOR_NOR2_NUM785 (.ZN (N2531), .A1 (N2395), .A2 (N2458));
      NOR2_X1 XNOR_NOR2_NUM786 (.ZN (N2532), .A1 (N2458), .A2 (N1083));
      NOR2_X1 XNOR_NOR2_NUM787 (.ZN (N2533), .A1 (N2313), .A2 (N2458));
      NOR2_X1 XNOR_NOR2_NUM788 (.ZN (N2536), .A1 (N2462), .A2 (N2463));
      NOR2_X1 XNOR_NOR2_NUM789 (.ZN (N2539), .A1 (N2467), .A2 (N2464));
      NOR2_X1 XNOR_NOR2_NUM790 (.ZN (N2543), .A1 (N2407), .A2 (N2470));
      NOR2_X1 XNOR_NOR2_NUM791 (.ZN (N2544), .A1 (N2470), .A2 (N2404));
      NOR2_X1 XNOR_NOR2_NUM792 (.ZN (N2545), .A1 (N2474), .A2 (N2475));
      NOR2_X1 XNOR_NOR2_NUM793 (.ZN (N2548), .A1 (N2476), .A2 (N2477));
      NOR2_X1 XNOR_NOR2_NUM794 (.ZN (N2549), .A1 (N2481), .A2 (N2482));
      NOR2_X1 XNOR_NOR2_NUM795 (.ZN (N2552), .A1 (N2486), .A2 (N2487));
      NOR2_X1 XNOR_NOR2_NUM796 (.ZN (N2555), .A1 (N2491), .A2 (N2492));
      NOR2_X1 XNOR_NOR2_NUM797 (.ZN (N2558), .A1 (N2496), .A2 (N2497));
      NOR2_X1 XNOR_NOR2_NUM798 (.ZN (N2561), .A1 (N2501), .A2 (N2502));
      NOR2_X1 XNOR_NOR2_NUM799 (.ZN (N2564), .A1 (N2506), .A2 (N2507));
      NOR2_X1 XNOR_NOR2_NUM800 (.ZN (N2567), .A1 (N2511), .A2 (N2512));
      NOR2_X1 XNOR_NOR2_NUM801 (.ZN (N2570), .A1 (N2516), .A2 (N2517));
      NOR2_X1 XNOR_NOR2_NUM802 (.ZN (N2573), .A1 (N2521), .A2 (N2522));
      NOR2_X1 XNOR_NOR2_NUM803 (.ZN (N2576), .A1 (N2526), .A2 (N2527));
      NOR2_X1 XNOR_NOR2_NUM804 (.ZN (N2579), .A1 (N2531), .A2 (N2532));
      NOR2_X1 XNOR_NOR2_NUM805 (.ZN (N2582), .A1 (N2536), .A2 (N2533));
      NOR2_X1 XNOR_NOR2_NUM806 (.ZN (N2586), .A1 (N2467), .A2 (N2539));
      NOR2_X1 XNOR_NOR2_NUM807 (.ZN (N2587), .A1 (N2539), .A2 (N2464));
      NOR2_X1 XNOR_NOR2_NUM808 (.ZN (N2588), .A1 (N2543), .A2 (N2544));
      NOR2_X1 XNOR_NOR2_NUM809 (.ZN (N2591), .A1 (N2545), .A2 (N1230));
      NOR2_X1 XNOR_NOR2_NUM810 (.ZN (N2595), .A1 (N2549), .A2 (N2478));
      NOR2_X1 XNOR_NOR2_NUM811 (.ZN (N2599), .A1 (N2552), .A2 (N2483));
      NOR2_X1 XNOR_NOR2_NUM812 (.ZN (N2603), .A1 (N2555), .A2 (N2488));
      NOR2_X1 XNOR_NOR2_NUM813 (.ZN (N2607), .A1 (N2558), .A2 (N2493));
      NOR2_X1 XNOR_NOR2_NUM814 (.ZN (N2611), .A1 (N2561), .A2 (N2498));
      NOR2_X1 XNOR_NOR2_NUM815 (.ZN (N2615), .A1 (N2564), .A2 (N2503));
      NOR2_X1 XNOR_NOR2_NUM816 (.ZN (N2619), .A1 (N2567), .A2 (N2508));
      NOR2_X1 XNOR_NOR2_NUM817 (.ZN (N2623), .A1 (N2570), .A2 (N2513));
      NOR2_X1 XNOR_NOR2_NUM818 (.ZN (N2627), .A1 (N2573), .A2 (N2518));
      NOR2_X1 XNOR_NOR2_NUM819 (.ZN (N2631), .A1 (N2576), .A2 (N2523));
      NOR2_X1 XNOR_NOR2_NUM820 (.ZN (N2635), .A1 (N2579), .A2 (N2528));
      NOR2_X1 XNOR_NOR2_NUM821 (.ZN (N2639), .A1 (N2536), .A2 (N2582));
      NOR2_X1 XNOR_NOR2_NUM822 (.ZN (N2640), .A1 (N2582), .A2 (N2533));
      NOR2_X1 XNOR_NOR2_NUM823 (.ZN (N2641), .A1 (N2586), .A2 (N2587));
      NOR2_X1 XNOR_NOR2_NUM824 (.ZN (N2644), .A1 (N2588), .A2 (N1182));
      NOR2_X1 XNOR_NOR2_NUM825 (.ZN (N2648), .A1 (N2545), .A2 (N2591));
      NOR2_X1 XNOR_NOR2_NUM826 (.ZN (N2649), .A1 (N2591), .A2 (N1230));
      NOR2_X1 XNOR_NOR2_NUM827 (.ZN (N2650), .A1 (N2410), .A2 (N2591));
      NOR2_X1 XNOR_NOR2_NUM828 (.ZN (N2653), .A1 (N2549), .A2 (N2595));
      NOR2_X1 XNOR_NOR2_NUM829 (.ZN (N2654), .A1 (N2595), .A2 (N2478));
      NOR2_X1 XNOR_NOR2_NUM830 (.ZN (N2655), .A1 (N2552), .A2 (N2599));
      NOR2_X1 XNOR_NOR2_NUM831 (.ZN (N2656), .A1 (N2599), .A2 (N2483));
      NOR2_X1 XNOR_NOR2_NUM832 (.ZN (N2657), .A1 (N2555), .A2 (N2603));
      NOR2_X1 XNOR_NOR2_NUM833 (.ZN (N2658), .A1 (N2603), .A2 (N2488));
      NOR2_X1 XNOR_NOR2_NUM834 (.ZN (N2659), .A1 (N2558), .A2 (N2607));
      NOR2_X1 XNOR_NOR2_NUM835 (.ZN (N2660), .A1 (N2607), .A2 (N2493));
      NOR2_X1 XNOR_NOR2_NUM836 (.ZN (N2661), .A1 (N2561), .A2 (N2611));
      NOR2_X1 XNOR_NOR2_NUM837 (.ZN (N2662), .A1 (N2611), .A2 (N2498));
      NOR2_X1 XNOR_NOR2_NUM838 (.ZN (N2663), .A1 (N2564), .A2 (N2615));
      NOR2_X1 XNOR_NOR2_NUM839 (.ZN (N2664), .A1 (N2615), .A2 (N2503));
      NOR2_X1 XNOR_NOR2_NUM840 (.ZN (N2665), .A1 (N2567), .A2 (N2619));
      NOR2_X1 XNOR_NOR2_NUM841 (.ZN (N2666), .A1 (N2619), .A2 (N2508));
      NOR2_X1 XNOR_NOR2_NUM842 (.ZN (N2667), .A1 (N2570), .A2 (N2623));
      NOR2_X1 XNOR_NOR2_NUM843 (.ZN (N2668), .A1 (N2623), .A2 (N2513));
      NOR2_X1 XNOR_NOR2_NUM844 (.ZN (N2669), .A1 (N2573), .A2 (N2627));
      NOR2_X1 XNOR_NOR2_NUM845 (.ZN (N2670), .A1 (N2627), .A2 (N2518));
      NOR2_X1 XNOR_NOR2_NUM846 (.ZN (N2671), .A1 (N2576), .A2 (N2631));
      NOR2_X1 XNOR_NOR2_NUM847 (.ZN (N2672), .A1 (N2631), .A2 (N2523));
      NOR2_X1 XNOR_NOR2_NUM848 (.ZN (N2673), .A1 (N2579), .A2 (N2635));
      NOR2_X1 XNOR_NOR2_NUM849 (.ZN (N2674), .A1 (N2635), .A2 (N2528));
      NOR2_X1 XNOR_NOR2_NUM850 (.ZN (N2675), .A1 (N2639), .A2 (N2640));
      NOR2_X1 XNOR_NOR2_NUM851 (.ZN (N2678), .A1 (N2641), .A2 (N1134));
      NOR2_X1 XNOR_NOR2_NUM852 (.ZN (N2682), .A1 (N2588), .A2 (N2644));
      NOR2_X1 XNOR_NOR2_NUM853 (.ZN (N2683), .A1 (N2644), .A2 (N1182));
      NOR2_X1 XNOR_NOR2_NUM854 (.ZN (N2684), .A1 (N2470), .A2 (N2644));
      NOR2_X1 XNOR_NOR2_NUM855 (.ZN (N2687), .A1 (N2648), .A2 (N2649));
      NOR2_X1 XNOR_NOR2_NUM856 (.ZN (N2690), .A1 (N1278), .A2 (N2650));
      NOR2_X1 XNOR_NOR2_NUM857 (.ZN (N2694), .A1 (N2653), .A2 (N2654));
      NOR2_X1 XNOR_NOR2_NUM858 (.ZN (N2697), .A1 (N2655), .A2 (N2656));
      NOR2_X1 XNOR_NOR2_NUM859 (.ZN (N2700), .A1 (N2657), .A2 (N2658));
      NOR2_X1 XNOR_NOR2_NUM860 (.ZN (N2703), .A1 (N2659), .A2 (N2660));
      NOR2_X1 XNOR_NOR2_NUM861 (.ZN (N2706), .A1 (N2661), .A2 (N2662));
      NOR2_X1 XNOR_NOR2_NUM862 (.ZN (N2709), .A1 (N2663), .A2 (N2664));
      NOR2_X1 XNOR_NOR2_NUM863 (.ZN (N2712), .A1 (N2665), .A2 (N2666));
      NOR2_X1 XNOR_NOR2_NUM864 (.ZN (N2715), .A1 (N2667), .A2 (N2668));
      NOR2_X1 XNOR_NOR2_NUM865 (.ZN (N2718), .A1 (N2669), .A2 (N2670));
      NOR2_X1 XNOR_NOR2_NUM866 (.ZN (N2721), .A1 (N2671), .A2 (N2672));
      NOR2_X1 XNOR_NOR2_NUM867 (.ZN (N2724), .A1 (N2673), .A2 (N2674));
      NOR2_X1 XNOR_NOR2_NUM868 (.ZN (N2727), .A1 (N2675), .A2 (N1086));
      NOR2_X1 XNOR_NOR2_NUM869 (.ZN (N2731), .A1 (N2641), .A2 (N2678));
      NOR2_X1 XNOR_NOR2_NUM870 (.ZN (N2732), .A1 (N2678), .A2 (N1134));
      NOR2_X1 XNOR_NOR2_NUM871 (.ZN (N2733), .A1 (N2539), .A2 (N2678));
      NOR2_X1 XNOR_NOR2_NUM872 (.ZN (N2736), .A1 (N2682), .A2 (N2683));
      NOR2_X1 XNOR_NOR2_NUM873 (.ZN (N2739), .A1 (N2687), .A2 (N2684));
      NOR2_X1 XNOR_NOR2_NUM874 (.ZN (N2743), .A1 (N1278), .A2 (N2690));
      NOR2_X1 XNOR_NOR2_NUM875 (.ZN (N2744), .A1 (N2690), .A2 (N2650));
      NOR2_X1 XNOR_NOR2_NUM876 (.ZN (N2745), .A1 (N2694), .A2 (N558));
      NOR2_X1 XNOR_NOR2_NUM877 (.ZN (N2749), .A1 (N2697), .A2 (N606));
      NOR2_X1 XNOR_NOR2_NUM878 (.ZN (N2753), .A1 (N2700), .A2 (N654));
      NOR2_X1 XNOR_NOR2_NUM879 (.ZN (N2757), .A1 (N2703), .A2 (N702));
      NOR2_X1 XNOR_NOR2_NUM880 (.ZN (N2761), .A1 (N2706), .A2 (N750));
      NOR2_X1 XNOR_NOR2_NUM881 (.ZN (N2765), .A1 (N2709), .A2 (N798));
      NOR2_X1 XNOR_NOR2_NUM882 (.ZN (N2769), .A1 (N2712), .A2 (N846));
      NOR2_X1 XNOR_NOR2_NUM883 (.ZN (N2773), .A1 (N2715), .A2 (N894));
      NOR2_X1 XNOR_NOR2_NUM884 (.ZN (N2777), .A1 (N2718), .A2 (N942));
      NOR2_X1 XNOR_NOR2_NUM885 (.ZN (N2781), .A1 (N2721), .A2 (N990));
      NOR2_X1 XNOR_NOR2_NUM886 (.ZN (N2785), .A1 (N2724), .A2 (N1038));
      NOR2_X1 XNOR_NOR2_NUM887 (.ZN (N2789), .A1 (N2675), .A2 (N2727));
      NOR2_X1 XNOR_NOR2_NUM888 (.ZN (N2790), .A1 (N2727), .A2 (N1086));
      NOR2_X1 XNOR_NOR2_NUM889 (.ZN (N2791), .A1 (N2582), .A2 (N2727));
      NOR2_X1 XNOR_NOR2_NUM890 (.ZN (N2794), .A1 (N2731), .A2 (N2732));
      NOR2_X1 XNOR_NOR2_NUM891 (.ZN (N2797), .A1 (N2736), .A2 (N2733));
      NOR2_X1 XNOR_NOR2_NUM892 (.ZN (N2801), .A1 (N2687), .A2 (N2739));
      NOR2_X1 XNOR_NOR2_NUM893 (.ZN (N2802), .A1 (N2739), .A2 (N2684));
      NOR2_X1 XNOR_NOR2_NUM894 (.ZN (N2803), .A1 (N2743), .A2 (N2744));
      NOR2_X1 XNOR_NOR2_NUM895 (.ZN (N2806), .A1 (N2694), .A2 (N2745));
      NOR2_X1 XNOR_NOR2_NUM896 (.ZN (N2807), .A1 (N2745), .A2 (N558));
      NOR2_X1 XNOR_NOR2_NUM897 (.ZN (N2808), .A1 (N2595), .A2 (N2745));
      NOR2_X1 XNOR_NOR2_NUM898 (.ZN (N2811), .A1 (N2697), .A2 (N2749));
      NOR2_X1 XNOR_NOR2_NUM899 (.ZN (N2812), .A1 (N2749), .A2 (N606));
      NOR2_X1 XNOR_NOR2_NUM900 (.ZN (N2813), .A1 (N2599), .A2 (N2749));
      NOR2_X1 XNOR_NOR2_NUM901 (.ZN (N2816), .A1 (N2700), .A2 (N2753));
      NOR2_X1 XNOR_NOR2_NUM902 (.ZN (N2817), .A1 (N2753), .A2 (N654));
      NOR2_X1 XNOR_NOR2_NUM903 (.ZN (N2818), .A1 (N2603), .A2 (N2753));
      NOR2_X1 XNOR_NOR2_NUM904 (.ZN (N2821), .A1 (N2703), .A2 (N2757));
      NOR2_X1 XNOR_NOR2_NUM905 (.ZN (N2822), .A1 (N2757), .A2 (N702));
      NOR2_X1 XNOR_NOR2_NUM906 (.ZN (N2823), .A1 (N2607), .A2 (N2757));
      NOR2_X1 XNOR_NOR2_NUM907 (.ZN (N2826), .A1 (N2706), .A2 (N2761));
      NOR2_X1 XNOR_NOR2_NUM908 (.ZN (N2827), .A1 (N2761), .A2 (N750));
      NOR2_X1 XNOR_NOR2_NUM909 (.ZN (N2828), .A1 (N2611), .A2 (N2761));
      NOR2_X1 XNOR_NOR2_NUM910 (.ZN (N2831), .A1 (N2709), .A2 (N2765));
      NOR2_X1 XNOR_NOR2_NUM911 (.ZN (N2832), .A1 (N2765), .A2 (N798));
      NOR2_X1 XNOR_NOR2_NUM912 (.ZN (N2833), .A1 (N2615), .A2 (N2765));
      NOR2_X1 XNOR_NOR2_NUM913 (.ZN (N2836), .A1 (N2712), .A2 (N2769));
      NOR2_X1 XNOR_NOR2_NUM914 (.ZN (N2837), .A1 (N2769), .A2 (N846));
      NOR2_X1 XNOR_NOR2_NUM915 (.ZN (N2838), .A1 (N2619), .A2 (N2769));
      NOR2_X1 XNOR_NOR2_NUM916 (.ZN (N2841), .A1 (N2715), .A2 (N2773));
      NOR2_X1 XNOR_NOR2_NUM917 (.ZN (N2842), .A1 (N2773), .A2 (N894));
      NOR2_X1 XNOR_NOR2_NUM918 (.ZN (N2843), .A1 (N2623), .A2 (N2773));
      NOR2_X1 XNOR_NOR2_NUM919 (.ZN (N2846), .A1 (N2718), .A2 (N2777));
      NOR2_X1 XNOR_NOR2_NUM920 (.ZN (N2847), .A1 (N2777), .A2 (N942));
      NOR2_X1 XNOR_NOR2_NUM921 (.ZN (N2848), .A1 (N2627), .A2 (N2777));
      NOR2_X1 XNOR_NOR2_NUM922 (.ZN (N2851), .A1 (N2721), .A2 (N2781));
      NOR2_X1 XNOR_NOR2_NUM923 (.ZN (N2852), .A1 (N2781), .A2 (N990));
      NOR2_X1 XNOR_NOR2_NUM924 (.ZN (N2853), .A1 (N2631), .A2 (N2781));
      NOR2_X1 XNOR_NOR2_NUM925 (.ZN (N2856), .A1 (N2724), .A2 (N2785));
      NOR2_X1 XNOR_NOR2_NUM926 (.ZN (N2857), .A1 (N2785), .A2 (N1038));
      NOR2_X1 XNOR_NOR2_NUM927 (.ZN (N2858), .A1 (N2635), .A2 (N2785));
      NOR2_X1 XNOR_NOR2_NUM928 (.ZN (N2861), .A1 (N2789), .A2 (N2790));
      NOR2_X1 XNOR_NOR2_NUM929 (.ZN (N2864), .A1 (N2794), .A2 (N2791));
      NOR2_X1 XNOR_NOR2_NUM930 (.ZN (N2868), .A1 (N2736), .A2 (N2797));
      NOR2_X1 XNOR_NOR2_NUM931 (.ZN (N2869), .A1 (N2797), .A2 (N2733));
      NOR2_X1 XNOR_NOR2_NUM932 (.ZN (N2870), .A1 (N2801), .A2 (N2802));
      NOR2_X1 XNOR_NOR2_NUM933 (.ZN (N2873), .A1 (N2803), .A2 (N1233));
      NOR2_X1 XNOR_NOR2_NUM934 (.ZN (N2877), .A1 (N2806), .A2 (N2807));
      NOR2_X1 XNOR_NOR2_NUM935 (.ZN (N2878), .A1 (N2811), .A2 (N2812));
      NOR2_X1 XNOR_NOR2_NUM936 (.ZN (N2881), .A1 (N2816), .A2 (N2817));
      NOR2_X1 XNOR_NOR2_NUM937 (.ZN (N2884), .A1 (N2821), .A2 (N2822));
      NOR2_X1 XNOR_NOR2_NUM938 (.ZN (N2887), .A1 (N2826), .A2 (N2827));
      NOR2_X1 XNOR_NOR2_NUM939 (.ZN (N2890), .A1 (N2831), .A2 (N2832));
      NOR2_X1 XNOR_NOR2_NUM940 (.ZN (N2893), .A1 (N2836), .A2 (N2837));
      NOR2_X1 XNOR_NOR2_NUM941 (.ZN (N2896), .A1 (N2841), .A2 (N2842));
      NOR2_X1 XNOR_NOR2_NUM942 (.ZN (N2899), .A1 (N2846), .A2 (N2847));
      NOR2_X1 XNOR_NOR2_NUM943 (.ZN (N2902), .A1 (N2851), .A2 (N2852));
      NOR2_X1 XNOR_NOR2_NUM944 (.ZN (N2905), .A1 (N2856), .A2 (N2857));
      NOR2_X1 XNOR_NOR2_NUM945 (.ZN (N2908), .A1 (N2861), .A2 (N2858));
      NOR2_X1 XNOR_NOR2_NUM946 (.ZN (N2912), .A1 (N2794), .A2 (N2864));
      NOR2_X1 XNOR_NOR2_NUM947 (.ZN (N2913), .A1 (N2864), .A2 (N2791));
      NOR2_X1 XNOR_NOR2_NUM948 (.ZN (N2914), .A1 (N2868), .A2 (N2869));
      NOR2_X1 XNOR_NOR2_NUM949 (.ZN (N2917), .A1 (N2870), .A2 (N1185));
      NOR2_X1 XNOR_NOR2_NUM950 (.ZN (N2921), .A1 (N2803), .A2 (N2873));
      NOR2_X1 XNOR_NOR2_NUM951 (.ZN (N2922), .A1 (N2873), .A2 (N1233));
      NOR2_X1 XNOR_NOR2_NUM952 (.ZN (N2923), .A1 (N2690), .A2 (N2873));
      NOR2_X1 XNOR_NOR2_NUM953 (.ZN (N2926), .A1 (N2878), .A2 (N2808));
      NOR2_X1 XNOR_NOR2_NUM954 (.ZN (N2930), .A1 (N2881), .A2 (N2813));
      NOR2_X1 XNOR_NOR2_NUM955 (.ZN (N2934), .A1 (N2884), .A2 (N2818));
      NOR2_X1 XNOR_NOR2_NUM956 (.ZN (N2938), .A1 (N2887), .A2 (N2823));
      NOR2_X1 XNOR_NOR2_NUM957 (.ZN (N2942), .A1 (N2890), .A2 (N2828));
      NOR2_X1 XNOR_NOR2_NUM958 (.ZN (N2946), .A1 (N2893), .A2 (N2833));
      NOR2_X1 XNOR_NOR2_NUM959 (.ZN (N2950), .A1 (N2896), .A2 (N2838));
      NOR2_X1 XNOR_NOR2_NUM960 (.ZN (N2954), .A1 (N2899), .A2 (N2843));
      NOR2_X1 XNOR_NOR2_NUM961 (.ZN (N2958), .A1 (N2902), .A2 (N2848));
      NOR2_X1 XNOR_NOR2_NUM962 (.ZN (N2962), .A1 (N2905), .A2 (N2853));
      NOR2_X1 XNOR_NOR2_NUM963 (.ZN (N2966), .A1 (N2861), .A2 (N2908));
      NOR2_X1 XNOR_NOR2_NUM964 (.ZN (N2967), .A1 (N2908), .A2 (N2858));
      NOR2_X1 XNOR_NOR2_NUM965 (.ZN (N2968), .A1 (N2912), .A2 (N2913));
      NOR2_X1 XNOR_NOR2_NUM966 (.ZN (N2971), .A1 (N2914), .A2 (N1137));
      NOR2_X1 XNOR_NOR2_NUM967 (.ZN (N2975), .A1 (N2870), .A2 (N2917));
      NOR2_X1 XNOR_NOR2_NUM968 (.ZN (N2976), .A1 (N2917), .A2 (N1185));
      NOR2_X1 XNOR_NOR2_NUM969 (.ZN (N2977), .A1 (N2739), .A2 (N2917));
      NOR2_X1 XNOR_NOR2_NUM970 (.ZN (N2980), .A1 (N2921), .A2 (N2922));
      NOR2_X1 XNOR_NOR2_NUM971 (.ZN (N2983), .A1 (N1281), .A2 (N2923));
      NOR2_X1 XNOR_NOR2_NUM972 (.ZN (N2987), .A1 (N2878), .A2 (N2926));
      NOR2_X1 XNOR_NOR2_NUM973 (.ZN (N2988), .A1 (N2926), .A2 (N2808));
      NOR2_X1 XNOR_NOR2_NUM974 (.ZN (N2989), .A1 (N2881), .A2 (N2930));
      NOR2_X1 XNOR_NOR2_NUM975 (.ZN (N2990), .A1 (N2930), .A2 (N2813));
      NOR2_X1 XNOR_NOR2_NUM976 (.ZN (N2991), .A1 (N2884), .A2 (N2934));
      NOR2_X1 XNOR_NOR2_NUM977 (.ZN (N2992), .A1 (N2934), .A2 (N2818));
      NOR2_X1 XNOR_NOR2_NUM978 (.ZN (N2993), .A1 (N2887), .A2 (N2938));
      NOR2_X1 XNOR_NOR2_NUM979 (.ZN (N2994), .A1 (N2938), .A2 (N2823));
      NOR2_X1 XNOR_NOR2_NUM980 (.ZN (N2995), .A1 (N2890), .A2 (N2942));
      NOR2_X1 XNOR_NOR2_NUM981 (.ZN (N2996), .A1 (N2942), .A2 (N2828));
      NOR2_X1 XNOR_NOR2_NUM982 (.ZN (N2997), .A1 (N2893), .A2 (N2946));
      NOR2_X1 XNOR_NOR2_NUM983 (.ZN (N2998), .A1 (N2946), .A2 (N2833));
      NOR2_X1 XNOR_NOR2_NUM984 (.ZN (N2999), .A1 (N2896), .A2 (N2950));
      NOR2_X1 XNOR_NOR2_NUM985 (.ZN (N3000), .A1 (N2950), .A2 (N2838));
      NOR2_X1 XNOR_NOR2_NUM986 (.ZN (N3001), .A1 (N2899), .A2 (N2954));
      NOR2_X1 XNOR_NOR2_NUM987 (.ZN (N3002), .A1 (N2954), .A2 (N2843));
      NOR2_X1 XNOR_NOR2_NUM988 (.ZN (N3003), .A1 (N2902), .A2 (N2958));
      NOR2_X1 XNOR_NOR2_NUM989 (.ZN (N3004), .A1 (N2958), .A2 (N2848));
      NOR2_X1 XNOR_NOR2_NUM990 (.ZN (N3005), .A1 (N2905), .A2 (N2962));
      NOR2_X1 XNOR_NOR2_NUM991 (.ZN (N3006), .A1 (N2962), .A2 (N2853));
      NOR2_X1 XNOR_NOR2_NUM992 (.ZN (N3007), .A1 (N2966), .A2 (N2967));
      NOR2_X1 XNOR_NOR2_NUM993 (.ZN (N3010), .A1 (N2968), .A2 (N1089));
      NOR2_X1 XNOR_NOR2_NUM994 (.ZN (N3014), .A1 (N2914), .A2 (N2971));
      NOR2_X1 XNOR_NOR2_NUM995 (.ZN (N3015), .A1 (N2971), .A2 (N1137));
      NOR2_X1 XNOR_NOR2_NUM996 (.ZN (N3016), .A1 (N2797), .A2 (N2971));
      NOR2_X1 XNOR_NOR2_NUM997 (.ZN (N3019), .A1 (N2975), .A2 (N2976));
      NOR2_X1 XNOR_NOR2_NUM998 (.ZN (N3022), .A1 (N2980), .A2 (N2977));
      NOR2_X1 XNOR_NOR2_NUM999 (.ZN (N3026), .A1 (N1281), .A2 (N2983));
      NOR2_X1 XNOR_NOR2_NUM1000 (.ZN (N3027), .A1 (N2983), .A2 (N2923));
      NOR2_X1 XNOR_NOR2_NUM1001 (.ZN (N3028), .A1 (N2987), .A2 (N2988));
      NOR2_X1 XNOR_NOR2_NUM1002 (.ZN (N3031), .A1 (N2989), .A2 (N2990));
      NOR2_X1 XNOR_NOR2_NUM1003 (.ZN (N3034), .A1 (N2991), .A2 (N2992));
      NOR2_X1 XNOR_NOR2_NUM1004 (.ZN (N3037), .A1 (N2993), .A2 (N2994));
      NOR2_X1 XNOR_NOR2_NUM1005 (.ZN (N3040), .A1 (N2995), .A2 (N2996));
      NOR2_X1 XNOR_NOR2_NUM1006 (.ZN (N3043), .A1 (N2997), .A2 (N2998));
      NOR2_X1 XNOR_NOR2_NUM1007 (.ZN (N3046), .A1 (N2999), .A2 (N3000));
      NOR2_X1 XNOR_NOR2_NUM1008 (.ZN (N3049), .A1 (N3001), .A2 (N3002));
      NOR2_X1 XNOR_NOR2_NUM1009 (.ZN (N3052), .A1 (N3003), .A2 (N3004));
      NOR2_X1 XNOR_NOR2_NUM1010 (.ZN (N3055), .A1 (N3005), .A2 (N3006));
      NOR2_X1 XNOR_NOR2_NUM1011 (.ZN (N3058), .A1 (N3007), .A2 (N1041));
      NOR2_X1 XNOR_NOR2_NUM1012 (.ZN (N3062), .A1 (N2968), .A2 (N3010));
      NOR2_X1 XNOR_NOR2_NUM1013 (.ZN (N3063), .A1 (N3010), .A2 (N1089));
      NOR2_X1 XNOR_NOR2_NUM1014 (.ZN (N3064), .A1 (N2864), .A2 (N3010));
      NOR2_X1 XNOR_NOR2_NUM1015 (.ZN (N3067), .A1 (N3014), .A2 (N3015));
      NOR2_X1 XNOR_NOR2_NUM1016 (.ZN (N3070), .A1 (N3019), .A2 (N3016));
      NOR2_X1 XNOR_NOR2_NUM1017 (.ZN (N3074), .A1 (N2980), .A2 (N3022));
      NOR2_X1 XNOR_NOR2_NUM1018 (.ZN (N3075), .A1 (N3022), .A2 (N2977));
      NOR2_X1 XNOR_NOR2_NUM1019 (.ZN (N3076), .A1 (N3026), .A2 (N3027));
      NOR2_X1 XNOR_NOR2_NUM1020 (.ZN (N3079), .A1 (N3028), .A2 (N561));
      NOR2_X1 XNOR_NOR2_NUM1021 (.ZN (N3083), .A1 (N3031), .A2 (N609));
      NOR2_X1 XNOR_NOR2_NUM1022 (.ZN (N3087), .A1 (N3034), .A2 (N657));
      NOR2_X1 XNOR_NOR2_NUM1023 (.ZN (N3091), .A1 (N3037), .A2 (N705));
      NOR2_X1 XNOR_NOR2_NUM1024 (.ZN (N3095), .A1 (N3040), .A2 (N753));
      NOR2_X1 XNOR_NOR2_NUM1025 (.ZN (N3099), .A1 (N3043), .A2 (N801));
      NOR2_X1 XNOR_NOR2_NUM1026 (.ZN (N3103), .A1 (N3046), .A2 (N849));
      NOR2_X1 XNOR_NOR2_NUM1027 (.ZN (N3107), .A1 (N3049), .A2 (N897));
      NOR2_X1 XNOR_NOR2_NUM1028 (.ZN (N3111), .A1 (N3052), .A2 (N945));
      NOR2_X1 XNOR_NOR2_NUM1029 (.ZN (N3115), .A1 (N3055), .A2 (N993));
      NOR2_X1 XNOR_NOR2_NUM1030 (.ZN (N3119), .A1 (N3007), .A2 (N3058));
      NOR2_X1 XNOR_NOR2_NUM1031 (.ZN (N3120), .A1 (N3058), .A2 (N1041));
      NOR2_X1 XNOR_NOR2_NUM1032 (.ZN (N3121), .A1 (N2908), .A2 (N3058));
      NOR2_X1 XNOR_NOR2_NUM1033 (.ZN (N3124), .A1 (N3062), .A2 (N3063));
      NOR2_X1 XNOR_NOR2_NUM1034 (.ZN (N3127), .A1 (N3067), .A2 (N3064));
      NOR2_X1 XNOR_NOR2_NUM1035 (.ZN (N3131), .A1 (N3019), .A2 (N3070));
      NOR2_X1 XNOR_NOR2_NUM1036 (.ZN (N3132), .A1 (N3070), .A2 (N3016));
      NOR2_X1 XNOR_NOR2_NUM1037 (.ZN (N3133), .A1 (N3074), .A2 (N3075));
      NOR2_X1 XNOR_NOR2_NUM1038 (.ZN (N3136), .A1 (N3076), .A2 (N1236));
      NOR2_X1 XNOR_NOR2_NUM1039 (.ZN (N3140), .A1 (N3028), .A2 (N3079));
      NOR2_X1 XNOR_NOR2_NUM1040 (.ZN (N3141), .A1 (N3079), .A2 (N561));
      NOR2_X1 XNOR_NOR2_NUM1041 (.ZN (N3142), .A1 (N2926), .A2 (N3079));
      NOR2_X1 XNOR_NOR2_NUM1042 (.ZN (N3145), .A1 (N3031), .A2 (N3083));
      NOR2_X1 XNOR_NOR2_NUM1043 (.ZN (N3146), .A1 (N3083), .A2 (N609));
      NOR2_X1 XNOR_NOR2_NUM1044 (.ZN (N3147), .A1 (N2930), .A2 (N3083));
      NOR2_X1 XNOR_NOR2_NUM1045 (.ZN (N3150), .A1 (N3034), .A2 (N3087));
      NOR2_X1 XNOR_NOR2_NUM1046 (.ZN (N3151), .A1 (N3087), .A2 (N657));
      NOR2_X1 XNOR_NOR2_NUM1047 (.ZN (N3152), .A1 (N2934), .A2 (N3087));
      NOR2_X1 XNOR_NOR2_NUM1048 (.ZN (N3155), .A1 (N3037), .A2 (N3091));
      NOR2_X1 XNOR_NOR2_NUM1049 (.ZN (N3156), .A1 (N3091), .A2 (N705));
      NOR2_X1 XNOR_NOR2_NUM1050 (.ZN (N3157), .A1 (N2938), .A2 (N3091));
      NOR2_X1 XNOR_NOR2_NUM1051 (.ZN (N3160), .A1 (N3040), .A2 (N3095));
      NOR2_X1 XNOR_NOR2_NUM1052 (.ZN (N3161), .A1 (N3095), .A2 (N753));
      NOR2_X1 XNOR_NOR2_NUM1053 (.ZN (N3162), .A1 (N2942), .A2 (N3095));
      NOR2_X1 XNOR_NOR2_NUM1054 (.ZN (N3165), .A1 (N3043), .A2 (N3099));
      NOR2_X1 XNOR_NOR2_NUM1055 (.ZN (N3166), .A1 (N3099), .A2 (N801));
      NOR2_X1 XNOR_NOR2_NUM1056 (.ZN (N3167), .A1 (N2946), .A2 (N3099));
      NOR2_X1 XNOR_NOR2_NUM1057 (.ZN (N3170), .A1 (N3046), .A2 (N3103));
      NOR2_X1 XNOR_NOR2_NUM1058 (.ZN (N3171), .A1 (N3103), .A2 (N849));
      NOR2_X1 XNOR_NOR2_NUM1059 (.ZN (N3172), .A1 (N2950), .A2 (N3103));
      NOR2_X1 XNOR_NOR2_NUM1060 (.ZN (N3175), .A1 (N3049), .A2 (N3107));
      NOR2_X1 XNOR_NOR2_NUM1061 (.ZN (N3176), .A1 (N3107), .A2 (N897));
      NOR2_X1 XNOR_NOR2_NUM1062 (.ZN (N3177), .A1 (N2954), .A2 (N3107));
      NOR2_X1 XNOR_NOR2_NUM1063 (.ZN (N3180), .A1 (N3052), .A2 (N3111));
      NOR2_X1 XNOR_NOR2_NUM1064 (.ZN (N3181), .A1 (N3111), .A2 (N945));
      NOR2_X1 XNOR_NOR2_NUM1065 (.ZN (N3182), .A1 (N2958), .A2 (N3111));
      NOR2_X1 XNOR_NOR2_NUM1066 (.ZN (N3185), .A1 (N3055), .A2 (N3115));
      NOR2_X1 XNOR_NOR2_NUM1067 (.ZN (N3186), .A1 (N3115), .A2 (N993));
      NOR2_X1 XNOR_NOR2_NUM1068 (.ZN (N3187), .A1 (N2962), .A2 (N3115));
      NOR2_X1 XNOR_NOR2_NUM1069 (.ZN (N3190), .A1 (N3119), .A2 (N3120));
      NOR2_X1 XNOR_NOR2_NUM1070 (.ZN (N3193), .A1 (N3124), .A2 (N3121));
      NOR2_X1 XNOR_NOR2_NUM1071 (.ZN (N3197), .A1 (N3067), .A2 (N3127));
      NOR2_X1 XNOR_NOR2_NUM1072 (.ZN (N3198), .A1 (N3127), .A2 (N3064));
      NOR2_X1 XNOR_NOR2_NUM1073 (.ZN (N3199), .A1 (N3131), .A2 (N3132));
      NOR2_X1 XNOR_NOR2_NUM1074 (.ZN (N3202), .A1 (N3133), .A2 (N1188));
      NOR2_X1 XNOR_NOR2_NUM1075 (.ZN (N3206), .A1 (N3076), .A2 (N3136));
      NOR2_X1 XNOR_NOR2_NUM1076 (.ZN (N3207), .A1 (N3136), .A2 (N1236));
      NOR2_X1 XNOR_NOR2_NUM1077 (.ZN (N3208), .A1 (N2983), .A2 (N3136));
      NOR2_X1 XNOR_NOR2_NUM1078 (.ZN (N3211), .A1 (N3140), .A2 (N3141));
      NOR2_X1 XNOR_NOR2_NUM1079 (.ZN (N3212), .A1 (N3145), .A2 (N3146));
      NOR2_X1 XNOR_NOR2_NUM1080 (.ZN (N3215), .A1 (N3150), .A2 (N3151));
      NOR2_X1 XNOR_NOR2_NUM1081 (.ZN (N3218), .A1 (N3155), .A2 (N3156));
      NOR2_X1 XNOR_NOR2_NUM1082 (.ZN (N3221), .A1 (N3160), .A2 (N3161));
      NOR2_X1 XNOR_NOR2_NUM1083 (.ZN (N3224), .A1 (N3165), .A2 (N3166));
      NOR2_X1 XNOR_NOR2_NUM1084 (.ZN (N3227), .A1 (N3170), .A2 (N3171));
      NOR2_X1 XNOR_NOR2_NUM1085 (.ZN (N3230), .A1 (N3175), .A2 (N3176));
      NOR2_X1 XNOR_NOR2_NUM1086 (.ZN (N3233), .A1 (N3180), .A2 (N3181));
      NOR2_X1 XNOR_NOR2_NUM1087 (.ZN (N3236), .A1 (N3185), .A2 (N3186));
      NOR2_X1 XNOR_NOR2_NUM1088 (.ZN (N3239), .A1 (N3190), .A2 (N3187));
      NOR2_X1 XNOR_NOR2_NUM1089 (.ZN (N3243), .A1 (N3124), .A2 (N3193));
      NOR2_X1 XNOR_NOR2_NUM1090 (.ZN (N3244), .A1 (N3193), .A2 (N3121));
      NOR2_X1 XNOR_NOR2_NUM1091 (.ZN (N3245), .A1 (N3197), .A2 (N3198));
      NOR2_X1 XNOR_NOR2_NUM1092 (.ZN (N3248), .A1 (N3199), .A2 (N1140));
      NOR2_X1 XNOR_NOR2_NUM1093 (.ZN (N3252), .A1 (N3133), .A2 (N3202));
      NOR2_X1 XNOR_NOR2_NUM1094 (.ZN (N3253), .A1 (N3202), .A2 (N1188));
      NOR2_X1 XNOR_NOR2_NUM1095 (.ZN (N3254), .A1 (N3022), .A2 (N3202));
      NOR2_X1 XNOR_NOR2_NUM1096 (.ZN (N3257), .A1 (N3206), .A2 (N3207));
      NOR2_X1 XNOR_NOR2_NUM1097 (.ZN (N3260), .A1 (N1284), .A2 (N3208));
      NOR2_X1 XNOR_NOR2_NUM1098 (.ZN (N3264), .A1 (N3212), .A2 (N3142));
      NOR2_X1 XNOR_NOR2_NUM1099 (.ZN (N3268), .A1 (N3215), .A2 (N3147));
      NOR2_X1 XNOR_NOR2_NUM1100 (.ZN (N3272), .A1 (N3218), .A2 (N3152));
      NOR2_X1 XNOR_NOR2_NUM1101 (.ZN (N3276), .A1 (N3221), .A2 (N3157));
      NOR2_X1 XNOR_NOR2_NUM1102 (.ZN (N3280), .A1 (N3224), .A2 (N3162));
      NOR2_X1 XNOR_NOR2_NUM1103 (.ZN (N3284), .A1 (N3227), .A2 (N3167));
      NOR2_X1 XNOR_NOR2_NUM1104 (.ZN (N3288), .A1 (N3230), .A2 (N3172));
      NOR2_X1 XNOR_NOR2_NUM1105 (.ZN (N3292), .A1 (N3233), .A2 (N3177));
      NOR2_X1 XNOR_NOR2_NUM1106 (.ZN (N3296), .A1 (N3236), .A2 (N3182));
      NOR2_X1 XNOR_NOR2_NUM1107 (.ZN (N3300), .A1 (N3190), .A2 (N3239));
      NOR2_X1 XNOR_NOR2_NUM1108 (.ZN (N3301), .A1 (N3239), .A2 (N3187));
      NOR2_X1 XNOR_NOR2_NUM1109 (.ZN (N3302), .A1 (N3243), .A2 (N3244));
      NOR2_X1 XNOR_NOR2_NUM1110 (.ZN (N3305), .A1 (N3245), .A2 (N1092));
      NOR2_X1 XNOR_NOR2_NUM1111 (.ZN (N3309), .A1 (N3199), .A2 (N3248));
      NOR2_X1 XNOR_NOR2_NUM1112 (.ZN (N3310), .A1 (N3248), .A2 (N1140));
      NOR2_X1 XNOR_NOR2_NUM1113 (.ZN (N3311), .A1 (N3070), .A2 (N3248));
      NOR2_X1 XNOR_NOR2_NUM1114 (.ZN (N3314), .A1 (N3252), .A2 (N3253));
      NOR2_X1 XNOR_NOR2_NUM1115 (.ZN (N3317), .A1 (N3257), .A2 (N3254));
      NOR2_X1 XNOR_NOR2_NUM1116 (.ZN (N3321), .A1 (N1284), .A2 (N3260));
      NOR2_X1 XNOR_NOR2_NUM1117 (.ZN (N3322), .A1 (N3260), .A2 (N3208));
      NOR2_X1 XNOR_NOR2_NUM1118 (.ZN (N3323), .A1 (N3212), .A2 (N3264));
      NOR2_X1 XNOR_NOR2_NUM1119 (.ZN (N3324), .A1 (N3264), .A2 (N3142));
      NOR2_X1 XNOR_NOR2_NUM1120 (.ZN (N3325), .A1 (N3215), .A2 (N3268));
      NOR2_X1 XNOR_NOR2_NUM1121 (.ZN (N3326), .A1 (N3268), .A2 (N3147));
      NOR2_X1 XNOR_NOR2_NUM1122 (.ZN (N3327), .A1 (N3218), .A2 (N3272));
      NOR2_X1 XNOR_NOR2_NUM1123 (.ZN (N3328), .A1 (N3272), .A2 (N3152));
      NOR2_X1 XNOR_NOR2_NUM1124 (.ZN (N3329), .A1 (N3221), .A2 (N3276));
      NOR2_X1 XNOR_NOR2_NUM1125 (.ZN (N3330), .A1 (N3276), .A2 (N3157));
      NOR2_X1 XNOR_NOR2_NUM1126 (.ZN (N3331), .A1 (N3224), .A2 (N3280));
      NOR2_X1 XNOR_NOR2_NUM1127 (.ZN (N3332), .A1 (N3280), .A2 (N3162));
      NOR2_X1 XNOR_NOR2_NUM1128 (.ZN (N3333), .A1 (N3227), .A2 (N3284));
      NOR2_X1 XNOR_NOR2_NUM1129 (.ZN (N3334), .A1 (N3284), .A2 (N3167));
      NOR2_X1 XNOR_NOR2_NUM1130 (.ZN (N3335), .A1 (N3230), .A2 (N3288));
      NOR2_X1 XNOR_NOR2_NUM1131 (.ZN (N3336), .A1 (N3288), .A2 (N3172));
      NOR2_X1 XNOR_NOR2_NUM1132 (.ZN (N3337), .A1 (N3233), .A2 (N3292));
      NOR2_X1 XNOR_NOR2_NUM1133 (.ZN (N3338), .A1 (N3292), .A2 (N3177));
      NOR2_X1 XNOR_NOR2_NUM1134 (.ZN (N3339), .A1 (N3236), .A2 (N3296));
      NOR2_X1 XNOR_NOR2_NUM1135 (.ZN (N3340), .A1 (N3296), .A2 (N3182));
      NOR2_X1 XNOR_NOR2_NUM1136 (.ZN (N3341), .A1 (N3300), .A2 (N3301));
      NOR2_X1 XNOR_NOR2_NUM1137 (.ZN (N3344), .A1 (N3302), .A2 (N1044));
      NOR2_X1 XNOR_NOR2_NUM1138 (.ZN (N3348), .A1 (N3245), .A2 (N3305));
      NOR2_X1 XNOR_NOR2_NUM1139 (.ZN (N3349), .A1 (N3305), .A2 (N1092));
      NOR2_X1 XNOR_NOR2_NUM1140 (.ZN (N3350), .A1 (N3127), .A2 (N3305));
      NOR2_X1 XNOR_NOR2_NUM1141 (.ZN (N3353), .A1 (N3309), .A2 (N3310));
      NOR2_X1 XNOR_NOR2_NUM1142 (.ZN (N3356), .A1 (N3314), .A2 (N3311));
      NOR2_X1 XNOR_NOR2_NUM1143 (.ZN (N3360), .A1 (N3257), .A2 (N3317));
      NOR2_X1 XNOR_NOR2_NUM1144 (.ZN (N3361), .A1 (N3317), .A2 (N3254));
      NOR2_X1 XNOR_NOR2_NUM1145 (.ZN (N3362), .A1 (N3321), .A2 (N3322));
      NOR2_X1 XNOR_NOR2_NUM1146 (.ZN (N3365), .A1 (N3323), .A2 (N3324));
      NOR2_X1 XNOR_NOR2_NUM1147 (.ZN (N3368), .A1 (N3325), .A2 (N3326));
      NOR2_X1 XNOR_NOR2_NUM1148 (.ZN (N3371), .A1 (N3327), .A2 (N3328));
      NOR2_X1 XNOR_NOR2_NUM1149 (.ZN (N3374), .A1 (N3329), .A2 (N3330));
      NOR2_X1 XNOR_NOR2_NUM1150 (.ZN (N3377), .A1 (N3331), .A2 (N3332));
      NOR2_X1 XNOR_NOR2_NUM1151 (.ZN (N3380), .A1 (N3333), .A2 (N3334));
      NOR2_X1 XNOR_NOR2_NUM1152 (.ZN (N3383), .A1 (N3335), .A2 (N3336));
      NOR2_X1 XNOR_NOR2_NUM1153 (.ZN (N3386), .A1 (N3337), .A2 (N3338));
      NOR2_X1 XNOR_NOR2_NUM1154 (.ZN (N3389), .A1 (N3339), .A2 (N3340));
      NOR2_X1 XNOR_NOR2_NUM1155 (.ZN (N3392), .A1 (N3341), .A2 (N996));
      NOR2_X1 XNOR_NOR2_NUM1156 (.ZN (N3396), .A1 (N3302), .A2 (N3344));
      NOR2_X1 XNOR_NOR2_NUM1157 (.ZN (N3397), .A1 (N3344), .A2 (N1044));
      NOR2_X1 XNOR_NOR2_NUM1158 (.ZN (N3398), .A1 (N3193), .A2 (N3344));
      NOR2_X1 XNOR_NOR2_NUM1159 (.ZN (N3401), .A1 (N3348), .A2 (N3349));
      NOR2_X1 XNOR_NOR2_NUM1160 (.ZN (N3404), .A1 (N3353), .A2 (N3350));
      NOR2_X1 XNOR_NOR2_NUM1161 (.ZN (N3408), .A1 (N3314), .A2 (N3356));
      NOR2_X1 XNOR_NOR2_NUM1162 (.ZN (N3409), .A1 (N3356), .A2 (N3311));
      NOR2_X1 XNOR_NOR2_NUM1163 (.ZN (N3410), .A1 (N3360), .A2 (N3361));
      NOR2_X1 XNOR_NOR2_NUM1164 (.ZN (N3413), .A1 (N3362), .A2 (N1239));
      NOR2_X1 XNOR_NOR2_NUM1165 (.ZN (N3417), .A1 (N3365), .A2 (N564));
      NOR2_X1 XNOR_NOR2_NUM1166 (.ZN (N3421), .A1 (N3368), .A2 (N612));
      NOR2_X1 XNOR_NOR2_NUM1167 (.ZN (N3425), .A1 (N3371), .A2 (N660));
      NOR2_X1 XNOR_NOR2_NUM1168 (.ZN (N3429), .A1 (N3374), .A2 (N708));
      NOR2_X1 XNOR_NOR2_NUM1169 (.ZN (N3433), .A1 (N3377), .A2 (N756));
      NOR2_X1 XNOR_NOR2_NUM1170 (.ZN (N3437), .A1 (N3380), .A2 (N804));
      NOR2_X1 XNOR_NOR2_NUM1171 (.ZN (N3441), .A1 (N3383), .A2 (N852));
      NOR2_X1 XNOR_NOR2_NUM1172 (.ZN (N3445), .A1 (N3386), .A2 (N900));
      NOR2_X1 XNOR_NOR2_NUM1173 (.ZN (N3449), .A1 (N3389), .A2 (N948));
      NOR2_X1 XNOR_NOR2_NUM1174 (.ZN (N3453), .A1 (N3341), .A2 (N3392));
      NOR2_X1 XNOR_NOR2_NUM1175 (.ZN (N3454), .A1 (N3392), .A2 (N996));
      NOR2_X1 XNOR_NOR2_NUM1176 (.ZN (N3455), .A1 (N3239), .A2 (N3392));
      NOR2_X1 XNOR_NOR2_NUM1177 (.ZN (N3458), .A1 (N3396), .A2 (N3397));
      NOR2_X1 XNOR_NOR2_NUM1178 (.ZN (N3461), .A1 (N3401), .A2 (N3398));
      NOR2_X1 XNOR_NOR2_NUM1179 (.ZN (N3465), .A1 (N3353), .A2 (N3404));
      NOR2_X1 XNOR_NOR2_NUM1180 (.ZN (N3466), .A1 (N3404), .A2 (N3350));
      NOR2_X1 XNOR_NOR2_NUM1181 (.ZN (N3467), .A1 (N3408), .A2 (N3409));
      NOR2_X1 XNOR_NOR2_NUM1182 (.ZN (N3470), .A1 (N3410), .A2 (N1191));
      NOR2_X1 XNOR_NOR2_NUM1183 (.ZN (N3474), .A1 (N3362), .A2 (N3413));
      NOR2_X1 XNOR_NOR2_NUM1184 (.ZN (N3475), .A1 (N3413), .A2 (N1239));
      NOR2_X1 XNOR_NOR2_NUM1185 (.ZN (N3476), .A1 (N3260), .A2 (N3413));
      NOR2_X1 XNOR_NOR2_NUM1186 (.ZN (N3479), .A1 (N3365), .A2 (N3417));
      NOR2_X1 XNOR_NOR2_NUM1187 (.ZN (N3480), .A1 (N3417), .A2 (N564));
      NOR2_X1 XNOR_NOR2_NUM1188 (.ZN (N3481), .A1 (N3264), .A2 (N3417));
      NOR2_X1 XNOR_NOR2_NUM1189 (.ZN (N3484), .A1 (N3368), .A2 (N3421));
      NOR2_X1 XNOR_NOR2_NUM1190 (.ZN (N3485), .A1 (N3421), .A2 (N612));
      NOR2_X1 XNOR_NOR2_NUM1191 (.ZN (N3486), .A1 (N3268), .A2 (N3421));
      NOR2_X1 XNOR_NOR2_NUM1192 (.ZN (N3489), .A1 (N3371), .A2 (N3425));
      NOR2_X1 XNOR_NOR2_NUM1193 (.ZN (N3490), .A1 (N3425), .A2 (N660));
      NOR2_X1 XNOR_NOR2_NUM1194 (.ZN (N3491), .A1 (N3272), .A2 (N3425));
      NOR2_X1 XNOR_NOR2_NUM1195 (.ZN (N3494), .A1 (N3374), .A2 (N3429));
      NOR2_X1 XNOR_NOR2_NUM1196 (.ZN (N3495), .A1 (N3429), .A2 (N708));
      NOR2_X1 XNOR_NOR2_NUM1197 (.ZN (N3496), .A1 (N3276), .A2 (N3429));
      NOR2_X1 XNOR_NOR2_NUM1198 (.ZN (N3499), .A1 (N3377), .A2 (N3433));
      NOR2_X1 XNOR_NOR2_NUM1199 (.ZN (N3500), .A1 (N3433), .A2 (N756));
      NOR2_X1 XNOR_NOR2_NUM1200 (.ZN (N3501), .A1 (N3280), .A2 (N3433));
      NOR2_X1 XNOR_NOR2_NUM1201 (.ZN (N3504), .A1 (N3380), .A2 (N3437));
      NOR2_X1 XNOR_NOR2_NUM1202 (.ZN (N3505), .A1 (N3437), .A2 (N804));
      NOR2_X1 XNOR_NOR2_NUM1203 (.ZN (N3506), .A1 (N3284), .A2 (N3437));
      NOR2_X1 XNOR_NOR2_NUM1204 (.ZN (N3509), .A1 (N3383), .A2 (N3441));
      NOR2_X1 XNOR_NOR2_NUM1205 (.ZN (N3510), .A1 (N3441), .A2 (N852));
      NOR2_X1 XNOR_NOR2_NUM1206 (.ZN (N3511), .A1 (N3288), .A2 (N3441));
      NOR2_X1 XNOR_NOR2_NUM1207 (.ZN (N3514), .A1 (N3386), .A2 (N3445));
      NOR2_X1 XNOR_NOR2_NUM1208 (.ZN (N3515), .A1 (N3445), .A2 (N900));
      NOR2_X1 XNOR_NOR2_NUM1209 (.ZN (N3516), .A1 (N3292), .A2 (N3445));
      NOR2_X1 XNOR_NOR2_NUM1210 (.ZN (N3519), .A1 (N3389), .A2 (N3449));
      NOR2_X1 XNOR_NOR2_NUM1211 (.ZN (N3520), .A1 (N3449), .A2 (N948));
      NOR2_X1 XNOR_NOR2_NUM1212 (.ZN (N3521), .A1 (N3296), .A2 (N3449));
      NOR2_X1 XNOR_NOR2_NUM1213 (.ZN (N3524), .A1 (N3453), .A2 (N3454));
      NOR2_X1 XNOR_NOR2_NUM1214 (.ZN (N3527), .A1 (N3458), .A2 (N3455));
      NOR2_X1 XNOR_NOR2_NUM1215 (.ZN (N3531), .A1 (N3401), .A2 (N3461));
      NOR2_X1 XNOR_NOR2_NUM1216 (.ZN (N3532), .A1 (N3461), .A2 (N3398));
      NOR2_X1 XNOR_NOR2_NUM1217 (.ZN (N3533), .A1 (N3465), .A2 (N3466));
      NOR2_X1 XNOR_NOR2_NUM1218 (.ZN (N3536), .A1 (N3467), .A2 (N1143));
      NOR2_X1 XNOR_NOR2_NUM1219 (.ZN (N3540), .A1 (N3410), .A2 (N3470));
      NOR2_X1 XNOR_NOR2_NUM1220 (.ZN (N3541), .A1 (N3470), .A2 (N1191));
      NOR2_X1 XNOR_NOR2_NUM1221 (.ZN (N3542), .A1 (N3317), .A2 (N3470));
      NOR2_X1 XNOR_NOR2_NUM1222 (.ZN (N3545), .A1 (N3474), .A2 (N3475));
      NOR2_X1 XNOR_NOR2_NUM1223 (.ZN (N3548), .A1 (N1287), .A2 (N3476));
      NOR2_X1 XNOR_NOR2_NUM1224 (.ZN (N3552), .A1 (N3479), .A2 (N3480));
      NOR2_X1 XNOR_NOR2_NUM1225 (.ZN (N3553), .A1 (N3484), .A2 (N3485));
      NOR2_X1 XNOR_NOR2_NUM1226 (.ZN (N3556), .A1 (N3489), .A2 (N3490));
      NOR2_X1 XNOR_NOR2_NUM1227 (.ZN (N3559), .A1 (N3494), .A2 (N3495));
      NOR2_X1 XNOR_NOR2_NUM1228 (.ZN (N3562), .A1 (N3499), .A2 (N3500));
      NOR2_X1 XNOR_NOR2_NUM1229 (.ZN (N3565), .A1 (N3504), .A2 (N3505));
      NOR2_X1 XNOR_NOR2_NUM1230 (.ZN (N3568), .A1 (N3509), .A2 (N3510));
      NOR2_X1 XNOR_NOR2_NUM1231 (.ZN (N3571), .A1 (N3514), .A2 (N3515));
      NOR2_X1 XNOR_NOR2_NUM1232 (.ZN (N3574), .A1 (N3519), .A2 (N3520));
      NOR2_X1 XNOR_NOR2_NUM1233 (.ZN (N3577), .A1 (N3524), .A2 (N3521));
      NOR2_X1 XNOR_NOR2_NUM1234 (.ZN (N3581), .A1 (N3458), .A2 (N3527));
      NOR2_X1 XNOR_NOR2_NUM1235 (.ZN (N3582), .A1 (N3527), .A2 (N3455));
      NOR2_X1 XNOR_NOR2_NUM1236 (.ZN (N3583), .A1 (N3531), .A2 (N3532));
      NOR2_X1 XNOR_NOR2_NUM1237 (.ZN (N3586), .A1 (N3533), .A2 (N1095));
      NOR2_X1 XNOR_NOR2_NUM1238 (.ZN (N3590), .A1 (N3467), .A2 (N3536));
      NOR2_X1 XNOR_NOR2_NUM1239 (.ZN (N3591), .A1 (N3536), .A2 (N1143));
      NOR2_X1 XNOR_NOR2_NUM1240 (.ZN (N3592), .A1 (N3356), .A2 (N3536));
      NOR2_X1 XNOR_NOR2_NUM1241 (.ZN (N3595), .A1 (N3540), .A2 (N3541));
      NOR2_X1 XNOR_NOR2_NUM1242 (.ZN (N3598), .A1 (N3545), .A2 (N3542));
      NOR2_X1 XNOR_NOR2_NUM1243 (.ZN (N3602), .A1 (N1287), .A2 (N3548));
      NOR2_X1 XNOR_NOR2_NUM1244 (.ZN (N3603), .A1 (N3548), .A2 (N3476));
      NOR2_X1 XNOR_NOR2_NUM1245 (.ZN (N3604), .A1 (N3553), .A2 (N3481));
      NOR2_X1 XNOR_NOR2_NUM1246 (.ZN (N3608), .A1 (N3556), .A2 (N3486));
      NOR2_X1 XNOR_NOR2_NUM1247 (.ZN (N3612), .A1 (N3559), .A2 (N3491));
      NOR2_X1 XNOR_NOR2_NUM1248 (.ZN (N3616), .A1 (N3562), .A2 (N3496));
      NOR2_X1 XNOR_NOR2_NUM1249 (.ZN (N3620), .A1 (N3565), .A2 (N3501));
      NOR2_X1 XNOR_NOR2_NUM1250 (.ZN (N3624), .A1 (N3568), .A2 (N3506));
      NOR2_X1 XNOR_NOR2_NUM1251 (.ZN (N3628), .A1 (N3571), .A2 (N3511));
      NOR2_X1 XNOR_NOR2_NUM1252 (.ZN (N3632), .A1 (N3574), .A2 (N3516));
      NOR2_X1 XNOR_NOR2_NUM1253 (.ZN (N3636), .A1 (N3524), .A2 (N3577));
      NOR2_X1 XNOR_NOR2_NUM1254 (.ZN (N3637), .A1 (N3577), .A2 (N3521));
      NOR2_X1 XNOR_NOR2_NUM1255 (.ZN (N3638), .A1 (N3581), .A2 (N3582));
      NOR2_X1 XNOR_NOR2_NUM1256 (.ZN (N3641), .A1 (N3583), .A2 (N1047));
      NOR2_X1 XNOR_NOR2_NUM1257 (.ZN (N3645), .A1 (N3533), .A2 (N3586));
      NOR2_X1 XNOR_NOR2_NUM1258 (.ZN (N3646), .A1 (N3586), .A2 (N1095));
      NOR2_X1 XNOR_NOR2_NUM1259 (.ZN (N3647), .A1 (N3404), .A2 (N3586));
      NOR2_X1 XNOR_NOR2_NUM1260 (.ZN (N3650), .A1 (N3590), .A2 (N3591));
      NOR2_X1 XNOR_NOR2_NUM1261 (.ZN (N3653), .A1 (N3595), .A2 (N3592));
      NOR2_X1 XNOR_NOR2_NUM1262 (.ZN (N3657), .A1 (N3545), .A2 (N3598));
      NOR2_X1 XNOR_NOR2_NUM1263 (.ZN (N3658), .A1 (N3598), .A2 (N3542));
      NOR2_X1 XNOR_NOR2_NUM1264 (.ZN (N3659), .A1 (N3602), .A2 (N3603));
      NOR2_X1 XNOR_NOR2_NUM1265 (.ZN (N3662), .A1 (N3553), .A2 (N3604));
      NOR2_X1 XNOR_NOR2_NUM1266 (.ZN (N3663), .A1 (N3604), .A2 (N3481));
      NOR2_X1 XNOR_NOR2_NUM1267 (.ZN (N3664), .A1 (N3556), .A2 (N3608));
      NOR2_X1 XNOR_NOR2_NUM1268 (.ZN (N3665), .A1 (N3608), .A2 (N3486));
      NOR2_X1 XNOR_NOR2_NUM1269 (.ZN (N3666), .A1 (N3559), .A2 (N3612));
      NOR2_X1 XNOR_NOR2_NUM1270 (.ZN (N3667), .A1 (N3612), .A2 (N3491));
      NOR2_X1 XNOR_NOR2_NUM1271 (.ZN (N3668), .A1 (N3562), .A2 (N3616));
      NOR2_X1 XNOR_NOR2_NUM1272 (.ZN (N3669), .A1 (N3616), .A2 (N3496));
      NOR2_X1 XNOR_NOR2_NUM1273 (.ZN (N3670), .A1 (N3565), .A2 (N3620));
      NOR2_X1 XNOR_NOR2_NUM1274 (.ZN (N3671), .A1 (N3620), .A2 (N3501));
      NOR2_X1 XNOR_NOR2_NUM1275 (.ZN (N3672), .A1 (N3568), .A2 (N3624));
      NOR2_X1 XNOR_NOR2_NUM1276 (.ZN (N3673), .A1 (N3624), .A2 (N3506));
      NOR2_X1 XNOR_NOR2_NUM1277 (.ZN (N3674), .A1 (N3571), .A2 (N3628));
      NOR2_X1 XNOR_NOR2_NUM1278 (.ZN (N3675), .A1 (N3628), .A2 (N3511));
      NOR2_X1 XNOR_NOR2_NUM1279 (.ZN (N3676), .A1 (N3574), .A2 (N3632));
      NOR2_X1 XNOR_NOR2_NUM1280 (.ZN (N3677), .A1 (N3632), .A2 (N3516));
      NOR2_X1 XNOR_NOR2_NUM1281 (.ZN (N3678), .A1 (N3636), .A2 (N3637));
      NOR2_X1 XNOR_NOR2_NUM1282 (.ZN (N3681), .A1 (N3638), .A2 (N999));
      NOR2_X1 XNOR_NOR2_NUM1283 (.ZN (N3685), .A1 (N3583), .A2 (N3641));
      NOR2_X1 XNOR_NOR2_NUM1284 (.ZN (N3686), .A1 (N3641), .A2 (N1047));
      NOR2_X1 XNOR_NOR2_NUM1285 (.ZN (N3687), .A1 (N3461), .A2 (N3641));
      NOR2_X1 XNOR_NOR2_NUM1286 (.ZN (N3690), .A1 (N3645), .A2 (N3646));
      NOR2_X1 XNOR_NOR2_NUM1287 (.ZN (N3693), .A1 (N3650), .A2 (N3647));
      NOR2_X1 XNOR_NOR2_NUM1288 (.ZN (N3697), .A1 (N3595), .A2 (N3653));
      NOR2_X1 XNOR_NOR2_NUM1289 (.ZN (N3698), .A1 (N3653), .A2 (N3592));
      NOR2_X1 XNOR_NOR2_NUM1290 (.ZN (N3699), .A1 (N3657), .A2 (N3658));
      NOR2_X1 XNOR_NOR2_NUM1291 (.ZN (N3702), .A1 (N3659), .A2 (N1242));
      NOR2_X1 XNOR_NOR2_NUM1292 (.ZN (N3706), .A1 (N3662), .A2 (N3663));
      NOR2_X1 XNOR_NOR2_NUM1293 (.ZN (N3709), .A1 (N3664), .A2 (N3665));
      NOR2_X1 XNOR_NOR2_NUM1294 (.ZN (N3712), .A1 (N3666), .A2 (N3667));
      NOR2_X1 XNOR_NOR2_NUM1295 (.ZN (N3715), .A1 (N3668), .A2 (N3669));
      NOR2_X1 XNOR_NOR2_NUM1296 (.ZN (N3718), .A1 (N3670), .A2 (N3671));
      NOR2_X1 XNOR_NOR2_NUM1297 (.ZN (N3721), .A1 (N3672), .A2 (N3673));
      NOR2_X1 XNOR_NOR2_NUM1298 (.ZN (N3724), .A1 (N3674), .A2 (N3675));
      NOR2_X1 XNOR_NOR2_NUM1299 (.ZN (N3727), .A1 (N3676), .A2 (N3677));
      NOR2_X1 XNOR_NOR2_NUM1300 (.ZN (N3730), .A1 (N3678), .A2 (N951));
      NOR2_X1 XNOR_NOR2_NUM1301 (.ZN (N3734), .A1 (N3638), .A2 (N3681));
      NOR2_X1 XNOR_NOR2_NUM1302 (.ZN (N3735), .A1 (N3681), .A2 (N999));
      NOR2_X1 XNOR_NOR2_NUM1303 (.ZN (N3736), .A1 (N3527), .A2 (N3681));
      NOR2_X1 XNOR_NOR2_NUM1304 (.ZN (N3739), .A1 (N3685), .A2 (N3686));
      NOR2_X1 XNOR_NOR2_NUM1305 (.ZN (N3742), .A1 (N3690), .A2 (N3687));
      NOR2_X1 XNOR_NOR2_NUM1306 (.ZN (N3746), .A1 (N3650), .A2 (N3693));
      NOR2_X1 XNOR_NOR2_NUM1307 (.ZN (N3747), .A1 (N3693), .A2 (N3647));
      NOR2_X1 XNOR_NOR2_NUM1308 (.ZN (N3748), .A1 (N3697), .A2 (N3698));
      NOR2_X1 XNOR_NOR2_NUM1309 (.ZN (N3751), .A1 (N3699), .A2 (N1194));
      NOR2_X1 XNOR_NOR2_NUM1310 (.ZN (N3755), .A1 (N3659), .A2 (N3702));
      NOR2_X1 XNOR_NOR2_NUM1311 (.ZN (N3756), .A1 (N3702), .A2 (N1242));
      NOR2_X1 XNOR_NOR2_NUM1312 (.ZN (N3757), .A1 (N3548), .A2 (N3702));
      NOR2_X1 XNOR_NOR2_NUM1313 (.ZN (N3760), .A1 (N3706), .A2 (N567));
      NOR2_X1 XNOR_NOR2_NUM1314 (.ZN (N3764), .A1 (N3709), .A2 (N615));
      NOR2_X1 XNOR_NOR2_NUM1315 (.ZN (N3768), .A1 (N3712), .A2 (N663));
      NOR2_X1 XNOR_NOR2_NUM1316 (.ZN (N3772), .A1 (N3715), .A2 (N711));
      NOR2_X1 XNOR_NOR2_NUM1317 (.ZN (N3776), .A1 (N3718), .A2 (N759));
      NOR2_X1 XNOR_NOR2_NUM1318 (.ZN (N3780), .A1 (N3721), .A2 (N807));
      NOR2_X1 XNOR_NOR2_NUM1319 (.ZN (N3784), .A1 (N3724), .A2 (N855));
      NOR2_X1 XNOR_NOR2_NUM1320 (.ZN (N3788), .A1 (N3727), .A2 (N903));
      NOR2_X1 XNOR_NOR2_NUM1321 (.ZN (N3792), .A1 (N3678), .A2 (N3730));
      NOR2_X1 XNOR_NOR2_NUM1322 (.ZN (N3793), .A1 (N3730), .A2 (N951));
      NOR2_X1 XNOR_NOR2_NUM1323 (.ZN (N3794), .A1 (N3577), .A2 (N3730));
      NOR2_X1 XNOR_NOR2_NUM1324 (.ZN (N3797), .A1 (N3734), .A2 (N3735));
      NOR2_X1 XNOR_NOR2_NUM1325 (.ZN (N3800), .A1 (N3739), .A2 (N3736));
      NOR2_X1 XNOR_NOR2_NUM1326 (.ZN (N3804), .A1 (N3690), .A2 (N3742));
      NOR2_X1 XNOR_NOR2_NUM1327 (.ZN (N3805), .A1 (N3742), .A2 (N3687));
      NOR2_X1 XNOR_NOR2_NUM1328 (.ZN (N3806), .A1 (N3746), .A2 (N3747));
      NOR2_X1 XNOR_NOR2_NUM1329 (.ZN (N3809), .A1 (N3748), .A2 (N1146));
      NOR2_X1 XNOR_NOR2_NUM1330 (.ZN (N3813), .A1 (N3699), .A2 (N3751));
      NOR2_X1 XNOR_NOR2_NUM1331 (.ZN (N3814), .A1 (N3751), .A2 (N1194));
      NOR2_X1 XNOR_NOR2_NUM1332 (.ZN (N3815), .A1 (N3598), .A2 (N3751));
      NOR2_X1 XNOR_NOR2_NUM1333 (.ZN (N3818), .A1 (N3755), .A2 (N3756));
      NOR2_X1 XNOR_NOR2_NUM1334 (.ZN (N3821), .A1 (N1290), .A2 (N3757));
      NOR2_X1 XNOR_NOR2_NUM1335 (.ZN (N3825), .A1 (N3706), .A2 (N3760));
      NOR2_X1 XNOR_NOR2_NUM1336 (.ZN (N3826), .A1 (N3760), .A2 (N567));
      NOR2_X1 XNOR_NOR2_NUM1337 (.ZN (N3827), .A1 (N3604), .A2 (N3760));
      NOR2_X1 XNOR_NOR2_NUM1338 (.ZN (N3830), .A1 (N3709), .A2 (N3764));
      NOR2_X1 XNOR_NOR2_NUM1339 (.ZN (N3831), .A1 (N3764), .A2 (N615));
      NOR2_X1 XNOR_NOR2_NUM1340 (.ZN (N3832), .A1 (N3608), .A2 (N3764));
      NOR2_X1 XNOR_NOR2_NUM1341 (.ZN (N3835), .A1 (N3712), .A2 (N3768));
      NOR2_X1 XNOR_NOR2_NUM1342 (.ZN (N3836), .A1 (N3768), .A2 (N663));
      NOR2_X1 XNOR_NOR2_NUM1343 (.ZN (N3837), .A1 (N3612), .A2 (N3768));
      NOR2_X1 XNOR_NOR2_NUM1344 (.ZN (N3840), .A1 (N3715), .A2 (N3772));
      NOR2_X1 XNOR_NOR2_NUM1345 (.ZN (N3841), .A1 (N3772), .A2 (N711));
      NOR2_X1 XNOR_NOR2_NUM1346 (.ZN (N3842), .A1 (N3616), .A2 (N3772));
      NOR2_X1 XNOR_NOR2_NUM1347 (.ZN (N3845), .A1 (N3718), .A2 (N3776));
      NOR2_X1 XNOR_NOR2_NUM1348 (.ZN (N3846), .A1 (N3776), .A2 (N759));
      NOR2_X1 XNOR_NOR2_NUM1349 (.ZN (N3847), .A1 (N3620), .A2 (N3776));
      NOR2_X1 XNOR_NOR2_NUM1350 (.ZN (N3850), .A1 (N3721), .A2 (N3780));
      NOR2_X1 XNOR_NOR2_NUM1351 (.ZN (N3851), .A1 (N3780), .A2 (N807));
      NOR2_X1 XNOR_NOR2_NUM1352 (.ZN (N3852), .A1 (N3624), .A2 (N3780));
      NOR2_X1 XNOR_NOR2_NUM1353 (.ZN (N3855), .A1 (N3724), .A2 (N3784));
      NOR2_X1 XNOR_NOR2_NUM1354 (.ZN (N3856), .A1 (N3784), .A2 (N855));
      NOR2_X1 XNOR_NOR2_NUM1355 (.ZN (N3857), .A1 (N3628), .A2 (N3784));
      NOR2_X1 XNOR_NOR2_NUM1356 (.ZN (N3860), .A1 (N3727), .A2 (N3788));
      NOR2_X1 XNOR_NOR2_NUM1357 (.ZN (N3861), .A1 (N3788), .A2 (N903));
      NOR2_X1 XNOR_NOR2_NUM1358 (.ZN (N3862), .A1 (N3632), .A2 (N3788));
      NOR2_X1 XNOR_NOR2_NUM1359 (.ZN (N3865), .A1 (N3792), .A2 (N3793));
      NOR2_X1 XNOR_NOR2_NUM1360 (.ZN (N3868), .A1 (N3797), .A2 (N3794));
      NOR2_X1 XNOR_NOR2_NUM1361 (.ZN (N3872), .A1 (N3739), .A2 (N3800));
      NOR2_X1 XNOR_NOR2_NUM1362 (.ZN (N3873), .A1 (N3800), .A2 (N3736));
      NOR2_X1 XNOR_NOR2_NUM1363 (.ZN (N3874), .A1 (N3804), .A2 (N3805));
      NOR2_X1 XNOR_NOR2_NUM1364 (.ZN (N3877), .A1 (N3806), .A2 (N1098));
      NOR2_X1 XNOR_NOR2_NUM1365 (.ZN (N3881), .A1 (N3748), .A2 (N3809));
      NOR2_X1 XNOR_NOR2_NUM1366 (.ZN (N3882), .A1 (N3809), .A2 (N1146));
      NOR2_X1 XNOR_NOR2_NUM1367 (.ZN (N3883), .A1 (N3653), .A2 (N3809));
      NOR2_X1 XNOR_NOR2_NUM1368 (.ZN (N3886), .A1 (N3813), .A2 (N3814));
      NOR2_X1 XNOR_NOR2_NUM1369 (.ZN (N3889), .A1 (N3818), .A2 (N3815));
      NOR2_X1 XNOR_NOR2_NUM1370 (.ZN (N3893), .A1 (N1290), .A2 (N3821));
      NOR2_X1 XNOR_NOR2_NUM1371 (.ZN (N3894), .A1 (N3821), .A2 (N3757));
      NOR2_X1 XNOR_NOR2_NUM1372 (.ZN (N3895), .A1 (N3825), .A2 (N3826));
      NOR2_X1 XNOR_NOR2_NUM1373 (.ZN (N3896), .A1 (N3830), .A2 (N3831));
      NOR2_X1 XNOR_NOR2_NUM1374 (.ZN (N3899), .A1 (N3835), .A2 (N3836));
      NOR2_X1 XNOR_NOR2_NUM1375 (.ZN (N3902), .A1 (N3840), .A2 (N3841));
      NOR2_X1 XNOR_NOR2_NUM1376 (.ZN (N3905), .A1 (N3845), .A2 (N3846));
      NOR2_X1 XNOR_NOR2_NUM1377 (.ZN (N3908), .A1 (N3850), .A2 (N3851));
      NOR2_X1 XNOR_NOR2_NUM1378 (.ZN (N3911), .A1 (N3855), .A2 (N3856));
      NOR2_X1 XNOR_NOR2_NUM1379 (.ZN (N3914), .A1 (N3860), .A2 (N3861));
      NOR2_X1 XNOR_NOR2_NUM1380 (.ZN (N3917), .A1 (N3865), .A2 (N3862));
      NOR2_X1 XNOR_NOR2_NUM1381 (.ZN (N3921), .A1 (N3797), .A2 (N3868));
      NOR2_X1 XNOR_NOR2_NUM1382 (.ZN (N3922), .A1 (N3868), .A2 (N3794));
      NOR2_X1 XNOR_NOR2_NUM1383 (.ZN (N3923), .A1 (N3872), .A2 (N3873));
      NOR2_X1 XNOR_NOR2_NUM1384 (.ZN (N3926), .A1 (N3874), .A2 (N1050));
      NOR2_X1 XNOR_NOR2_NUM1385 (.ZN (N3930), .A1 (N3806), .A2 (N3877));
      NOR2_X1 XNOR_NOR2_NUM1386 (.ZN (N3931), .A1 (N3877), .A2 (N1098));
      NOR2_X1 XNOR_NOR2_NUM1387 (.ZN (N3932), .A1 (N3693), .A2 (N3877));
      NOR2_X1 XNOR_NOR2_NUM1388 (.ZN (N3935), .A1 (N3881), .A2 (N3882));
      NOR2_X1 XNOR_NOR2_NUM1389 (.ZN (N3938), .A1 (N3886), .A2 (N3883));
      NOR2_X1 XNOR_NOR2_NUM1390 (.ZN (N3942), .A1 (N3818), .A2 (N3889));
      NOR2_X1 XNOR_NOR2_NUM1391 (.ZN (N3943), .A1 (N3889), .A2 (N3815));
      NOR2_X1 XNOR_NOR2_NUM1392 (.ZN (N3944), .A1 (N3893), .A2 (N3894));
      NOR2_X1 XNOR_NOR2_NUM1393 (.ZN (N3947), .A1 (N3896), .A2 (N3827));
      NOR2_X1 XNOR_NOR2_NUM1394 (.ZN (N3951), .A1 (N3899), .A2 (N3832));
      NOR2_X1 XNOR_NOR2_NUM1395 (.ZN (N3955), .A1 (N3902), .A2 (N3837));
      NOR2_X1 XNOR_NOR2_NUM1396 (.ZN (N3959), .A1 (N3905), .A2 (N3842));
      NOR2_X1 XNOR_NOR2_NUM1397 (.ZN (N3963), .A1 (N3908), .A2 (N3847));
      NOR2_X1 XNOR_NOR2_NUM1398 (.ZN (N3967), .A1 (N3911), .A2 (N3852));
      NOR2_X1 XNOR_NOR2_NUM1399 (.ZN (N3971), .A1 (N3914), .A2 (N3857));
      NOR2_X1 XNOR_NOR2_NUM1400 (.ZN (N3975), .A1 (N3865), .A2 (N3917));
      NOR2_X1 XNOR_NOR2_NUM1401 (.ZN (N3976), .A1 (N3917), .A2 (N3862));
      NOR2_X1 XNOR_NOR2_NUM1402 (.ZN (N3977), .A1 (N3921), .A2 (N3922));
      NOR2_X1 XNOR_NOR2_NUM1403 (.ZN (N3980), .A1 (N3923), .A2 (N1002));
      NOR2_X1 XNOR_NOR2_NUM1404 (.ZN (N3984), .A1 (N3874), .A2 (N3926));
      NOR2_X1 XNOR_NOR2_NUM1405 (.ZN (N3985), .A1 (N3926), .A2 (N1050));
      NOR2_X1 XNOR_NOR2_NUM1406 (.ZN (N3986), .A1 (N3742), .A2 (N3926));
      NOR2_X1 XNOR_NOR2_NUM1407 (.ZN (N3989), .A1 (N3930), .A2 (N3931));
      NOR2_X1 XNOR_NOR2_NUM1408 (.ZN (N3992), .A1 (N3935), .A2 (N3932));
      NOR2_X1 XNOR_NOR2_NUM1409 (.ZN (N3996), .A1 (N3886), .A2 (N3938));
      NOR2_X1 XNOR_NOR2_NUM1410 (.ZN (N3997), .A1 (N3938), .A2 (N3883));
      NOR2_X1 XNOR_NOR2_NUM1411 (.ZN (N3998), .A1 (N3942), .A2 (N3943));
      NOR2_X1 XNOR_NOR2_NUM1412 (.ZN (N4001), .A1 (N3944), .A2 (N1245));
      NOR2_X1 XNOR_NOR2_NUM1413 (.ZN (N4005), .A1 (N3896), .A2 (N3947));
      NOR2_X1 XNOR_NOR2_NUM1414 (.ZN (N4006), .A1 (N3947), .A2 (N3827));
      NOR2_X1 XNOR_NOR2_NUM1415 (.ZN (N4007), .A1 (N3899), .A2 (N3951));
      NOR2_X1 XNOR_NOR2_NUM1416 (.ZN (N4008), .A1 (N3951), .A2 (N3832));
      NOR2_X1 XNOR_NOR2_NUM1417 (.ZN (N4009), .A1 (N3902), .A2 (N3955));
      NOR2_X1 XNOR_NOR2_NUM1418 (.ZN (N4010), .A1 (N3955), .A2 (N3837));
      NOR2_X1 XNOR_NOR2_NUM1419 (.ZN (N4011), .A1 (N3905), .A2 (N3959));
      NOR2_X1 XNOR_NOR2_NUM1420 (.ZN (N4012), .A1 (N3959), .A2 (N3842));
      NOR2_X1 XNOR_NOR2_NUM1421 (.ZN (N4013), .A1 (N3908), .A2 (N3963));
      NOR2_X1 XNOR_NOR2_NUM1422 (.ZN (N4014), .A1 (N3963), .A2 (N3847));
      NOR2_X1 XNOR_NOR2_NUM1423 (.ZN (N4015), .A1 (N3911), .A2 (N3967));
      NOR2_X1 XNOR_NOR2_NUM1424 (.ZN (N4016), .A1 (N3967), .A2 (N3852));
      NOR2_X1 XNOR_NOR2_NUM1425 (.ZN (N4017), .A1 (N3914), .A2 (N3971));
      NOR2_X1 XNOR_NOR2_NUM1426 (.ZN (N4018), .A1 (N3971), .A2 (N3857));
      NOR2_X1 XNOR_NOR2_NUM1427 (.ZN (N4019), .A1 (N3975), .A2 (N3976));
      NOR2_X1 XNOR_NOR2_NUM1428 (.ZN (N4022), .A1 (N3977), .A2 (N954));
      NOR2_X1 XNOR_NOR2_NUM1429 (.ZN (N4026), .A1 (N3923), .A2 (N3980));
      NOR2_X1 XNOR_NOR2_NUM1430 (.ZN (N4027), .A1 (N3980), .A2 (N1002));
      NOR2_X1 XNOR_NOR2_NUM1431 (.ZN (N4028), .A1 (N3800), .A2 (N3980));
      NOR2_X1 XNOR_NOR2_NUM1432 (.ZN (N4031), .A1 (N3984), .A2 (N3985));
      NOR2_X1 XNOR_NOR2_NUM1433 (.ZN (N4034), .A1 (N3989), .A2 (N3986));
      NOR2_X1 XNOR_NOR2_NUM1434 (.ZN (N4038), .A1 (N3935), .A2 (N3992));
      NOR2_X1 XNOR_NOR2_NUM1435 (.ZN (N4039), .A1 (N3992), .A2 (N3932));
      NOR2_X1 XNOR_NOR2_NUM1436 (.ZN (N4040), .A1 (N3996), .A2 (N3997));
      NOR2_X1 XNOR_NOR2_NUM1437 (.ZN (N4043), .A1 (N3998), .A2 (N1197));
      NOR2_X1 XNOR_NOR2_NUM1438 (.ZN (N4047), .A1 (N3944), .A2 (N4001));
      NOR2_X1 XNOR_NOR2_NUM1439 (.ZN (N4048), .A1 (N4001), .A2 (N1245));
      NOR2_X1 XNOR_NOR2_NUM1440 (.ZN (N4049), .A1 (N3821), .A2 (N4001));
      NOR2_X1 XNOR_NOR2_NUM1441 (.ZN (N4052), .A1 (N4005), .A2 (N4006));
      NOR2_X1 XNOR_NOR2_NUM1442 (.ZN (N4055), .A1 (N4007), .A2 (N4008));
      NOR2_X1 XNOR_NOR2_NUM1443 (.ZN (N4058), .A1 (N4009), .A2 (N4010));
      NOR2_X1 XNOR_NOR2_NUM1444 (.ZN (N4061), .A1 (N4011), .A2 (N4012));
      NOR2_X1 XNOR_NOR2_NUM1445 (.ZN (N4064), .A1 (N4013), .A2 (N4014));
      NOR2_X1 XNOR_NOR2_NUM1446 (.ZN (N4067), .A1 (N4015), .A2 (N4016));
      NOR2_X1 XNOR_NOR2_NUM1447 (.ZN (N4070), .A1 (N4017), .A2 (N4018));
      NOR2_X1 XNOR_NOR2_NUM1448 (.ZN (N4073), .A1 (N4019), .A2 (N906));
      NOR2_X1 XNOR_NOR2_NUM1449 (.ZN (N4077), .A1 (N3977), .A2 (N4022));
      NOR2_X1 XNOR_NOR2_NUM1450 (.ZN (N4078), .A1 (N4022), .A2 (N954));
      NOR2_X1 XNOR_NOR2_NUM1451 (.ZN (N4079), .A1 (N3868), .A2 (N4022));
      NOR2_X1 XNOR_NOR2_NUM1452 (.ZN (N4082), .A1 (N4026), .A2 (N4027));
      NOR2_X1 XNOR_NOR2_NUM1453 (.ZN (N4085), .A1 (N4031), .A2 (N4028));
      NOR2_X1 XNOR_NOR2_NUM1454 (.ZN (N4089), .A1 (N3989), .A2 (N4034));
      NOR2_X1 XNOR_NOR2_NUM1455 (.ZN (N4090), .A1 (N4034), .A2 (N3986));
      NOR2_X1 XNOR_NOR2_NUM1456 (.ZN (N4091), .A1 (N4038), .A2 (N4039));
      NOR2_X1 XNOR_NOR2_NUM1457 (.ZN (N4094), .A1 (N4040), .A2 (N1149));
      NOR2_X1 XNOR_NOR2_NUM1458 (.ZN (N4098), .A1 (N3998), .A2 (N4043));
      NOR2_X1 XNOR_NOR2_NUM1459 (.ZN (N4099), .A1 (N4043), .A2 (N1197));
      NOR2_X1 XNOR_NOR2_NUM1460 (.ZN (N4100), .A1 (N3889), .A2 (N4043));
      NOR2_X1 XNOR_NOR2_NUM1461 (.ZN (N4103), .A1 (N4047), .A2 (N4048));
      NOR2_X1 XNOR_NOR2_NUM1462 (.ZN (N4106), .A1 (N1293), .A2 (N4049));
      NOR2_X1 XNOR_NOR2_NUM1463 (.ZN (N4110), .A1 (N4052), .A2 (N570));
      NOR2_X1 XNOR_NOR2_NUM1464 (.ZN (N4114), .A1 (N4055), .A2 (N618));
      NOR2_X1 XNOR_NOR2_NUM1465 (.ZN (N4118), .A1 (N4058), .A2 (N666));
      NOR2_X1 XNOR_NOR2_NUM1466 (.ZN (N4122), .A1 (N4061), .A2 (N714));
      NOR2_X1 XNOR_NOR2_NUM1467 (.ZN (N4126), .A1 (N4064), .A2 (N762));
      NOR2_X1 XNOR_NOR2_NUM1468 (.ZN (N4130), .A1 (N4067), .A2 (N810));
      NOR2_X1 XNOR_NOR2_NUM1469 (.ZN (N4134), .A1 (N4070), .A2 (N858));
      NOR2_X1 XNOR_NOR2_NUM1470 (.ZN (N4138), .A1 (N4019), .A2 (N4073));
      NOR2_X1 XNOR_NOR2_NUM1471 (.ZN (N4139), .A1 (N4073), .A2 (N906));
      NOR2_X1 XNOR_NOR2_NUM1472 (.ZN (N4140), .A1 (N3917), .A2 (N4073));
      NOR2_X1 XNOR_NOR2_NUM1473 (.ZN (N4143), .A1 (N4077), .A2 (N4078));
      NOR2_X1 XNOR_NOR2_NUM1474 (.ZN (N4146), .A1 (N4082), .A2 (N4079));
      NOR2_X1 XNOR_NOR2_NUM1475 (.ZN (N4150), .A1 (N4031), .A2 (N4085));
      NOR2_X1 XNOR_NOR2_NUM1476 (.ZN (N4151), .A1 (N4085), .A2 (N4028));
      NOR2_X1 XNOR_NOR2_NUM1477 (.ZN (N4152), .A1 (N4089), .A2 (N4090));
      NOR2_X1 XNOR_NOR2_NUM1478 (.ZN (N4155), .A1 (N4091), .A2 (N1101));
      NOR2_X1 XNOR_NOR2_NUM1479 (.ZN (N4159), .A1 (N4040), .A2 (N4094));
      NOR2_X1 XNOR_NOR2_NUM1480 (.ZN (N4160), .A1 (N4094), .A2 (N1149));
      NOR2_X1 XNOR_NOR2_NUM1481 (.ZN (N4161), .A1 (N3938), .A2 (N4094));
      NOR2_X1 XNOR_NOR2_NUM1482 (.ZN (N4164), .A1 (N4098), .A2 (N4099));
      NOR2_X1 XNOR_NOR2_NUM1483 (.ZN (N4167), .A1 (N4103), .A2 (N4100));
      NOR2_X1 XNOR_NOR2_NUM1484 (.ZN (N4171), .A1 (N1293), .A2 (N4106));
      NOR2_X1 XNOR_NOR2_NUM1485 (.ZN (N4172), .A1 (N4106), .A2 (N4049));
      NOR2_X1 XNOR_NOR2_NUM1486 (.ZN (N4173), .A1 (N4052), .A2 (N4110));
      NOR2_X1 XNOR_NOR2_NUM1487 (.ZN (N4174), .A1 (N4110), .A2 (N570));
      NOR2_X1 XNOR_NOR2_NUM1488 (.ZN (N4175), .A1 (N3947), .A2 (N4110));
      NOR2_X1 XNOR_NOR2_NUM1489 (.ZN (N4178), .A1 (N4055), .A2 (N4114));
      NOR2_X1 XNOR_NOR2_NUM1490 (.ZN (N4179), .A1 (N4114), .A2 (N618));
      NOR2_X1 XNOR_NOR2_NUM1491 (.ZN (N4180), .A1 (N3951), .A2 (N4114));
      NOR2_X1 XNOR_NOR2_NUM1492 (.ZN (N4183), .A1 (N4058), .A2 (N4118));
      NOR2_X1 XNOR_NOR2_NUM1493 (.ZN (N4184), .A1 (N4118), .A2 (N666));
      NOR2_X1 XNOR_NOR2_NUM1494 (.ZN (N4185), .A1 (N3955), .A2 (N4118));
      NOR2_X1 XNOR_NOR2_NUM1495 (.ZN (N4188), .A1 (N4061), .A2 (N4122));
      NOR2_X1 XNOR_NOR2_NUM1496 (.ZN (N4189), .A1 (N4122), .A2 (N714));
      NOR2_X1 XNOR_NOR2_NUM1497 (.ZN (N4190), .A1 (N3959), .A2 (N4122));
      NOR2_X1 XNOR_NOR2_NUM1498 (.ZN (N4193), .A1 (N4064), .A2 (N4126));
      NOR2_X1 XNOR_NOR2_NUM1499 (.ZN (N4194), .A1 (N4126), .A2 (N762));
      NOR2_X1 XNOR_NOR2_NUM1500 (.ZN (N4195), .A1 (N3963), .A2 (N4126));
      NOR2_X1 XNOR_NOR2_NUM1501 (.ZN (N4198), .A1 (N4067), .A2 (N4130));
      NOR2_X1 XNOR_NOR2_NUM1502 (.ZN (N4199), .A1 (N4130), .A2 (N810));
      NOR2_X1 XNOR_NOR2_NUM1503 (.ZN (N4200), .A1 (N3967), .A2 (N4130));
      NOR2_X1 XNOR_NOR2_NUM1504 (.ZN (N4203), .A1 (N4070), .A2 (N4134));
      NOR2_X1 XNOR_NOR2_NUM1505 (.ZN (N4204), .A1 (N4134), .A2 (N858));
      NOR2_X1 XNOR_NOR2_NUM1506 (.ZN (N4205), .A1 (N3971), .A2 (N4134));
      NOR2_X1 XNOR_NOR2_NUM1507 (.ZN (N4208), .A1 (N4138), .A2 (N4139));
      NOR2_X1 XNOR_NOR2_NUM1508 (.ZN (N4211), .A1 (N4143), .A2 (N4140));
      NOR2_X1 XNOR_NOR2_NUM1509 (.ZN (N4215), .A1 (N4082), .A2 (N4146));
      NOR2_X1 XNOR_NOR2_NUM1510 (.ZN (N4216), .A1 (N4146), .A2 (N4079));
      NOR2_X1 XNOR_NOR2_NUM1511 (.ZN (N4217), .A1 (N4150), .A2 (N4151));
      NOR2_X1 XNOR_NOR2_NUM1512 (.ZN (N4220), .A1 (N4152), .A2 (N1053));
      NOR2_X1 XNOR_NOR2_NUM1513 (.ZN (N4224), .A1 (N4091), .A2 (N4155));
      NOR2_X1 XNOR_NOR2_NUM1514 (.ZN (N4225), .A1 (N4155), .A2 (N1101));
      NOR2_X1 XNOR_NOR2_NUM1515 (.ZN (N4226), .A1 (N3992), .A2 (N4155));
      NOR2_X1 XNOR_NOR2_NUM1516 (.ZN (N4229), .A1 (N4159), .A2 (N4160));
      NOR2_X1 XNOR_NOR2_NUM1517 (.ZN (N4232), .A1 (N4164), .A2 (N4161));
      NOR2_X1 XNOR_NOR2_NUM1518 (.ZN (N4236), .A1 (N4103), .A2 (N4167));
      NOR2_X1 XNOR_NOR2_NUM1519 (.ZN (N4237), .A1 (N4167), .A2 (N4100));
      NOR2_X1 XNOR_NOR2_NUM1520 (.ZN (N4238), .A1 (N4171), .A2 (N4172));
      NOR2_X1 XNOR_NOR2_NUM1521 (.ZN (N4241), .A1 (N4173), .A2 (N4174));
      NOR2_X1 XNOR_NOR2_NUM1522 (.ZN (N4242), .A1 (N4178), .A2 (N4179));
      NOR2_X1 XNOR_NOR2_NUM1523 (.ZN (N4245), .A1 (N4183), .A2 (N4184));
      NOR2_X1 XNOR_NOR2_NUM1524 (.ZN (N4248), .A1 (N4188), .A2 (N4189));
      NOR2_X1 XNOR_NOR2_NUM1525 (.ZN (N4251), .A1 (N4193), .A2 (N4194));
      NOR2_X1 XNOR_NOR2_NUM1526 (.ZN (N4254), .A1 (N4198), .A2 (N4199));
      NOR2_X1 XNOR_NOR2_NUM1527 (.ZN (N4257), .A1 (N4203), .A2 (N4204));
      NOR2_X1 XNOR_NOR2_NUM1528 (.ZN (N4260), .A1 (N4208), .A2 (N4205));
      NOR2_X1 XNOR_NOR2_NUM1529 (.ZN (N4264), .A1 (N4143), .A2 (N4211));
      NOR2_X1 XNOR_NOR2_NUM1530 (.ZN (N4265), .A1 (N4211), .A2 (N4140));
      NOR2_X1 XNOR_NOR2_NUM1531 (.ZN (N4266), .A1 (N4215), .A2 (N4216));
      NOR2_X1 XNOR_NOR2_NUM1532 (.ZN (N4269), .A1 (N4217), .A2 (N1005));
      NOR2_X1 XNOR_NOR2_NUM1533 (.ZN (N4273), .A1 (N4152), .A2 (N4220));
      NOR2_X1 XNOR_NOR2_NUM1534 (.ZN (N4274), .A1 (N4220), .A2 (N1053));
      NOR2_X1 XNOR_NOR2_NUM1535 (.ZN (N4275), .A1 (N4034), .A2 (N4220));
      NOR2_X1 XNOR_NOR2_NUM1536 (.ZN (N4278), .A1 (N4224), .A2 (N4225));
      NOR2_X1 XNOR_NOR2_NUM1537 (.ZN (N4281), .A1 (N4229), .A2 (N4226));
      NOR2_X1 XNOR_NOR2_NUM1538 (.ZN (N4285), .A1 (N4164), .A2 (N4232));
      NOR2_X1 XNOR_NOR2_NUM1539 (.ZN (N4286), .A1 (N4232), .A2 (N4161));
      NOR2_X1 XNOR_NOR2_NUM1540 (.ZN (N4287), .A1 (N4236), .A2 (N4237));
      NOR2_X1 XNOR_NOR2_NUM1541 (.ZN (N4290), .A1 (N4238), .A2 (N1248));
      NOR2_X1 XNOR_NOR2_NUM1542 (.ZN (N4294), .A1 (N4242), .A2 (N4175));
      NOR2_X1 XNOR_NOR2_NUM1543 (.ZN (N4298), .A1 (N4245), .A2 (N4180));
      NOR2_X1 XNOR_NOR2_NUM1544 (.ZN (N4302), .A1 (N4248), .A2 (N4185));
      NOR2_X1 XNOR_NOR2_NUM1545 (.ZN (N4306), .A1 (N4251), .A2 (N4190));
      NOR2_X1 XNOR_NOR2_NUM1546 (.ZN (N4310), .A1 (N4254), .A2 (N4195));
      NOR2_X1 XNOR_NOR2_NUM1547 (.ZN (N4314), .A1 (N4257), .A2 (N4200));
      NOR2_X1 XNOR_NOR2_NUM1548 (.ZN (N4318), .A1 (N4208), .A2 (N4260));
      NOR2_X1 XNOR_NOR2_NUM1549 (.ZN (N4319), .A1 (N4260), .A2 (N4205));
      NOR2_X1 XNOR_NOR2_NUM1550 (.ZN (N4320), .A1 (N4264), .A2 (N4265));
      NOR2_X1 XNOR_NOR2_NUM1551 (.ZN (N4323), .A1 (N4266), .A2 (N957));
      NOR2_X1 XNOR_NOR2_NUM1552 (.ZN (N4327), .A1 (N4217), .A2 (N4269));
      NOR2_X1 XNOR_NOR2_NUM1553 (.ZN (N4328), .A1 (N4269), .A2 (N1005));
      NOR2_X1 XNOR_NOR2_NUM1554 (.ZN (N4329), .A1 (N4085), .A2 (N4269));
      NOR2_X1 XNOR_NOR2_NUM1555 (.ZN (N4332), .A1 (N4273), .A2 (N4274));
      NOR2_X1 XNOR_NOR2_NUM1556 (.ZN (N4335), .A1 (N4278), .A2 (N4275));
      NOR2_X1 XNOR_NOR2_NUM1557 (.ZN (N4339), .A1 (N4229), .A2 (N4281));
      NOR2_X1 XNOR_NOR2_NUM1558 (.ZN (N4340), .A1 (N4281), .A2 (N4226));
      NOR2_X1 XNOR_NOR2_NUM1559 (.ZN (N4341), .A1 (N4285), .A2 (N4286));
      NOR2_X1 XNOR_NOR2_NUM1560 (.ZN (N4344), .A1 (N4287), .A2 (N1200));
      NOR2_X1 XNOR_NOR2_NUM1561 (.ZN (N4348), .A1 (N4238), .A2 (N4290));
      NOR2_X1 XNOR_NOR2_NUM1562 (.ZN (N4349), .A1 (N4290), .A2 (N1248));
      NOR2_X1 XNOR_NOR2_NUM1563 (.ZN (N4350), .A1 (N4106), .A2 (N4290));
      NOR2_X1 XNOR_NOR2_NUM1564 (.ZN (N4353), .A1 (N4242), .A2 (N4294));
      NOR2_X1 XNOR_NOR2_NUM1565 (.ZN (N4354), .A1 (N4294), .A2 (N4175));
      NOR2_X1 XNOR_NOR2_NUM1566 (.ZN (N4355), .A1 (N4245), .A2 (N4298));
      NOR2_X1 XNOR_NOR2_NUM1567 (.ZN (N4356), .A1 (N4298), .A2 (N4180));
      NOR2_X1 XNOR_NOR2_NUM1568 (.ZN (N4357), .A1 (N4248), .A2 (N4302));
      NOR2_X1 XNOR_NOR2_NUM1569 (.ZN (N4358), .A1 (N4302), .A2 (N4185));
      NOR2_X1 XNOR_NOR2_NUM1570 (.ZN (N4359), .A1 (N4251), .A2 (N4306));
      NOR2_X1 XNOR_NOR2_NUM1571 (.ZN (N4360), .A1 (N4306), .A2 (N4190));
      NOR2_X1 XNOR_NOR2_NUM1572 (.ZN (N4361), .A1 (N4254), .A2 (N4310));
      NOR2_X1 XNOR_NOR2_NUM1573 (.ZN (N4362), .A1 (N4310), .A2 (N4195));
      NOR2_X1 XNOR_NOR2_NUM1574 (.ZN (N4363), .A1 (N4257), .A2 (N4314));
      NOR2_X1 XNOR_NOR2_NUM1575 (.ZN (N4364), .A1 (N4314), .A2 (N4200));
      NOR2_X1 XNOR_NOR2_NUM1576 (.ZN (N4365), .A1 (N4318), .A2 (N4319));
      NOR2_X1 XNOR_NOR2_NUM1577 (.ZN (N4368), .A1 (N4320), .A2 (N909));
      NOR2_X1 XNOR_NOR2_NUM1578 (.ZN (N4372), .A1 (N4266), .A2 (N4323));
      NOR2_X1 XNOR_NOR2_NUM1579 (.ZN (N4373), .A1 (N4323), .A2 (N957));
      NOR2_X1 XNOR_NOR2_NUM1580 (.ZN (N4374), .A1 (N4146), .A2 (N4323));
      NOR2_X1 XNOR_NOR2_NUM1581 (.ZN (N4377), .A1 (N4327), .A2 (N4328));
      NOR2_X1 XNOR_NOR2_NUM1582 (.ZN (N4380), .A1 (N4332), .A2 (N4329));
      NOR2_X1 XNOR_NOR2_NUM1583 (.ZN (N4384), .A1 (N4278), .A2 (N4335));
      NOR2_X1 XNOR_NOR2_NUM1584 (.ZN (N4385), .A1 (N4335), .A2 (N4275));
      NOR2_X1 XNOR_NOR2_NUM1585 (.ZN (N4386), .A1 (N4339), .A2 (N4340));
      NOR2_X1 XNOR_NOR2_NUM1586 (.ZN (N4389), .A1 (N4341), .A2 (N1152));
      NOR2_X1 XNOR_NOR2_NUM1587 (.ZN (N4393), .A1 (N4287), .A2 (N4344));
      NOR2_X1 XNOR_NOR2_NUM1588 (.ZN (N4394), .A1 (N4344), .A2 (N1200));
      NOR2_X1 XNOR_NOR2_NUM1589 (.ZN (N4395), .A1 (N4167), .A2 (N4344));
      NOR2_X1 XNOR_NOR2_NUM1590 (.ZN (N4398), .A1 (N4348), .A2 (N4349));
      NOR2_X1 XNOR_NOR2_NUM1591 (.ZN (N4401), .A1 (N1296), .A2 (N4350));
      NOR2_X1 XNOR_NOR2_NUM1592 (.ZN (N4405), .A1 (N4353), .A2 (N4354));
      NOR2_X1 XNOR_NOR2_NUM1593 (.ZN (N4408), .A1 (N4355), .A2 (N4356));
      NOR2_X1 XNOR_NOR2_NUM1594 (.ZN (N4411), .A1 (N4357), .A2 (N4358));
      NOR2_X1 XNOR_NOR2_NUM1595 (.ZN (N4414), .A1 (N4359), .A2 (N4360));
      NOR2_X1 XNOR_NOR2_NUM1596 (.ZN (N4417), .A1 (N4361), .A2 (N4362));
      NOR2_X1 XNOR_NOR2_NUM1597 (.ZN (N4420), .A1 (N4363), .A2 (N4364));
      NOR2_X1 XNOR_NOR2_NUM1598 (.ZN (N4423), .A1 (N4365), .A2 (N861));
      NOR2_X1 XNOR_NOR2_NUM1599 (.ZN (N4427), .A1 (N4320), .A2 (N4368));
      NOR2_X1 XNOR_NOR2_NUM1600 (.ZN (N4428), .A1 (N4368), .A2 (N909));
      NOR2_X1 XNOR_NOR2_NUM1601 (.ZN (N4429), .A1 (N4211), .A2 (N4368));
      NOR2_X1 XNOR_NOR2_NUM1602 (.ZN (N4432), .A1 (N4372), .A2 (N4373));
      NOR2_X1 XNOR_NOR2_NUM1603 (.ZN (N4435), .A1 (N4377), .A2 (N4374));
      NOR2_X1 XNOR_NOR2_NUM1604 (.ZN (N4439), .A1 (N4332), .A2 (N4380));
      NOR2_X1 XNOR_NOR2_NUM1605 (.ZN (N4440), .A1 (N4380), .A2 (N4329));
      NOR2_X1 XNOR_NOR2_NUM1606 (.ZN (N4441), .A1 (N4384), .A2 (N4385));
      NOR2_X1 XNOR_NOR2_NUM1607 (.ZN (N4444), .A1 (N4386), .A2 (N1104));
      NOR2_X1 XNOR_NOR2_NUM1608 (.ZN (N4448), .A1 (N4341), .A2 (N4389));
      NOR2_X1 XNOR_NOR2_NUM1609 (.ZN (N4449), .A1 (N4389), .A2 (N1152));
      NOR2_X1 XNOR_NOR2_NUM1610 (.ZN (N4450), .A1 (N4232), .A2 (N4389));
      NOR2_X1 XNOR_NOR2_NUM1611 (.ZN (N4453), .A1 (N4393), .A2 (N4394));
      NOR2_X1 XNOR_NOR2_NUM1612 (.ZN (N4456), .A1 (N4398), .A2 (N4395));
      NOR2_X1 XNOR_NOR2_NUM1613 (.ZN (N4460), .A1 (N1296), .A2 (N4401));
      NOR2_X1 XNOR_NOR2_NUM1614 (.ZN (N4461), .A1 (N4401), .A2 (N4350));
      NOR2_X1 XNOR_NOR2_NUM1615 (.ZN (N4462), .A1 (N4405), .A2 (N573));
      NOR2_X1 XNOR_NOR2_NUM1616 (.ZN (N4466), .A1 (N4408), .A2 (N621));
      NOR2_X1 XNOR_NOR2_NUM1617 (.ZN (N4470), .A1 (N4411), .A2 (N669));
      NOR2_X1 XNOR_NOR2_NUM1618 (.ZN (N4474), .A1 (N4414), .A2 (N717));
      NOR2_X1 XNOR_NOR2_NUM1619 (.ZN (N4478), .A1 (N4417), .A2 (N765));
      NOR2_X1 XNOR_NOR2_NUM1620 (.ZN (N4482), .A1 (N4420), .A2 (N813));
      NOR2_X1 XNOR_NOR2_NUM1621 (.ZN (N4486), .A1 (N4365), .A2 (N4423));
      NOR2_X1 XNOR_NOR2_NUM1622 (.ZN (N4487), .A1 (N4423), .A2 (N861));
      NOR2_X1 XNOR_NOR2_NUM1623 (.ZN (N4488), .A1 (N4260), .A2 (N4423));
      NOR2_X1 XNOR_NOR2_NUM1624 (.ZN (N4491), .A1 (N4427), .A2 (N4428));
      NOR2_X1 XNOR_NOR2_NUM1625 (.ZN (N4494), .A1 (N4432), .A2 (N4429));
      NOR2_X1 XNOR_NOR2_NUM1626 (.ZN (N4498), .A1 (N4377), .A2 (N4435));
      NOR2_X1 XNOR_NOR2_NUM1627 (.ZN (N4499), .A1 (N4435), .A2 (N4374));
      NOR2_X1 XNOR_NOR2_NUM1628 (.ZN (N4500), .A1 (N4439), .A2 (N4440));
      NOR2_X1 XNOR_NOR2_NUM1629 (.ZN (N4503), .A1 (N4441), .A2 (N1056));
      NOR2_X1 XNOR_NOR2_NUM1630 (.ZN (N4507), .A1 (N4386), .A2 (N4444));
      NOR2_X1 XNOR_NOR2_NUM1631 (.ZN (N4508), .A1 (N4444), .A2 (N1104));
      NOR2_X1 XNOR_NOR2_NUM1632 (.ZN (N4509), .A1 (N4281), .A2 (N4444));
      NOR2_X1 XNOR_NOR2_NUM1633 (.ZN (N4512), .A1 (N4448), .A2 (N4449));
      NOR2_X1 XNOR_NOR2_NUM1634 (.ZN (N4515), .A1 (N4453), .A2 (N4450));
      NOR2_X1 XNOR_NOR2_NUM1635 (.ZN (N4519), .A1 (N4398), .A2 (N4456));
      NOR2_X1 XNOR_NOR2_NUM1636 (.ZN (N4520), .A1 (N4456), .A2 (N4395));
      NOR2_X1 XNOR_NOR2_NUM1637 (.ZN (N4521), .A1 (N4460), .A2 (N4461));
      NOR2_X1 XNOR_NOR2_NUM1638 (.ZN (N4524), .A1 (N4405), .A2 (N4462));
      NOR2_X1 XNOR_NOR2_NUM1639 (.ZN (N4525), .A1 (N4462), .A2 (N573));
      NOR2_X1 XNOR_NOR2_NUM1640 (.ZN (N4526), .A1 (N4294), .A2 (N4462));
      NOR2_X1 XNOR_NOR2_NUM1641 (.ZN (N4529), .A1 (N4408), .A2 (N4466));
      NOR2_X1 XNOR_NOR2_NUM1642 (.ZN (N4530), .A1 (N4466), .A2 (N621));
      NOR2_X1 XNOR_NOR2_NUM1643 (.ZN (N4531), .A1 (N4298), .A2 (N4466));
      NOR2_X1 XNOR_NOR2_NUM1644 (.ZN (N4534), .A1 (N4411), .A2 (N4470));
      NOR2_X1 XNOR_NOR2_NUM1645 (.ZN (N4535), .A1 (N4470), .A2 (N669));
      NOR2_X1 XNOR_NOR2_NUM1646 (.ZN (N4536), .A1 (N4302), .A2 (N4470));
      NOR2_X1 XNOR_NOR2_NUM1647 (.ZN (N4539), .A1 (N4414), .A2 (N4474));
      NOR2_X1 XNOR_NOR2_NUM1648 (.ZN (N4540), .A1 (N4474), .A2 (N717));
      NOR2_X1 XNOR_NOR2_NUM1649 (.ZN (N4541), .A1 (N4306), .A2 (N4474));
      NOR2_X1 XNOR_NOR2_NUM1650 (.ZN (N4544), .A1 (N4417), .A2 (N4478));
      NOR2_X1 XNOR_NOR2_NUM1651 (.ZN (N4545), .A1 (N4478), .A2 (N765));
      NOR2_X1 XNOR_NOR2_NUM1652 (.ZN (N4546), .A1 (N4310), .A2 (N4478));
      NOR2_X1 XNOR_NOR2_NUM1653 (.ZN (N4549), .A1 (N4420), .A2 (N4482));
      NOR2_X1 XNOR_NOR2_NUM1654 (.ZN (N4550), .A1 (N4482), .A2 (N813));
      NOR2_X1 XNOR_NOR2_NUM1655 (.ZN (N4551), .A1 (N4314), .A2 (N4482));
      NOR2_X1 XNOR_NOR2_NUM1656 (.ZN (N4554), .A1 (N4486), .A2 (N4487));
      NOR2_X1 XNOR_NOR2_NUM1657 (.ZN (N4557), .A1 (N4491), .A2 (N4488));
      NOR2_X1 XNOR_NOR2_NUM1658 (.ZN (N4561), .A1 (N4432), .A2 (N4494));
      NOR2_X1 XNOR_NOR2_NUM1659 (.ZN (N4562), .A1 (N4494), .A2 (N4429));
      NOR2_X1 XNOR_NOR2_NUM1660 (.ZN (N4563), .A1 (N4498), .A2 (N4499));
      NOR2_X1 XNOR_NOR2_NUM1661 (.ZN (N4566), .A1 (N4500), .A2 (N1008));
      NOR2_X1 XNOR_NOR2_NUM1662 (.ZN (N4570), .A1 (N4441), .A2 (N4503));
      NOR2_X1 XNOR_NOR2_NUM1663 (.ZN (N4571), .A1 (N4503), .A2 (N1056));
      NOR2_X1 XNOR_NOR2_NUM1664 (.ZN (N4572), .A1 (N4335), .A2 (N4503));
      NOR2_X1 XNOR_NOR2_NUM1665 (.ZN (N4575), .A1 (N4507), .A2 (N4508));
      NOR2_X1 XNOR_NOR2_NUM1666 (.ZN (N4578), .A1 (N4512), .A2 (N4509));
      NOR2_X1 XNOR_NOR2_NUM1667 (.ZN (N4582), .A1 (N4453), .A2 (N4515));
      NOR2_X1 XNOR_NOR2_NUM1668 (.ZN (N4583), .A1 (N4515), .A2 (N4450));
      NOR2_X1 XNOR_NOR2_NUM1669 (.ZN (N4584), .A1 (N4519), .A2 (N4520));
      NOR2_X1 XNOR_NOR2_NUM1670 (.ZN (N4587), .A1 (N4521), .A2 (N1251));
      NOR2_X1 XNOR_NOR2_NUM1671 (.ZN (N4591), .A1 (N4524), .A2 (N4525));
      NOR2_X1 XNOR_NOR2_NUM1672 (.ZN (N4592), .A1 (N4529), .A2 (N4530));
      NOR2_X1 XNOR_NOR2_NUM1673 (.ZN (N4595), .A1 (N4534), .A2 (N4535));
      NOR2_X1 XNOR_NOR2_NUM1674 (.ZN (N4598), .A1 (N4539), .A2 (N4540));
      NOR2_X1 XNOR_NOR2_NUM1675 (.ZN (N4601), .A1 (N4544), .A2 (N4545));
      NOR2_X1 XNOR_NOR2_NUM1676 (.ZN (N4604), .A1 (N4549), .A2 (N4550));
      NOR2_X1 XNOR_NOR2_NUM1677 (.ZN (N4607), .A1 (N4554), .A2 (N4551));
      NOR2_X1 XNOR_NOR2_NUM1678 (.ZN (N4611), .A1 (N4491), .A2 (N4557));
      NOR2_X1 XNOR_NOR2_NUM1679 (.ZN (N4612), .A1 (N4557), .A2 (N4488));
      NOR2_X1 XNOR_NOR2_NUM1680 (.ZN (N4613), .A1 (N4561), .A2 (N4562));
      NOR2_X1 XNOR_NOR2_NUM1681 (.ZN (N4616), .A1 (N4563), .A2 (N960));
      NOR2_X1 XNOR_NOR2_NUM1682 (.ZN (N4620), .A1 (N4500), .A2 (N4566));
      NOR2_X1 XNOR_NOR2_NUM1683 (.ZN (N4621), .A1 (N4566), .A2 (N1008));
      NOR2_X1 XNOR_NOR2_NUM1684 (.ZN (N4622), .A1 (N4380), .A2 (N4566));
      NOR2_X1 XNOR_NOR2_NUM1685 (.ZN (N4625), .A1 (N4570), .A2 (N4571));
      NOR2_X1 XNOR_NOR2_NUM1686 (.ZN (N4628), .A1 (N4575), .A2 (N4572));
      NOR2_X1 XNOR_NOR2_NUM1687 (.ZN (N4632), .A1 (N4512), .A2 (N4578));
      NOR2_X1 XNOR_NOR2_NUM1688 (.ZN (N4633), .A1 (N4578), .A2 (N4509));
      NOR2_X1 XNOR_NOR2_NUM1689 (.ZN (N4634), .A1 (N4582), .A2 (N4583));
      NOR2_X1 XNOR_NOR2_NUM1690 (.ZN (N4637), .A1 (N4584), .A2 (N1203));
      NOR2_X1 XNOR_NOR2_NUM1691 (.ZN (N4641), .A1 (N4521), .A2 (N4587));
      NOR2_X1 XNOR_NOR2_NUM1692 (.ZN (N4642), .A1 (N4587), .A2 (N1251));
      NOR2_X1 XNOR_NOR2_NUM1693 (.ZN (N4643), .A1 (N4401), .A2 (N4587));
      NOR2_X1 XNOR_NOR2_NUM1694 (.ZN (N4646), .A1 (N4592), .A2 (N4526));
      NOR2_X1 XNOR_NOR2_NUM1695 (.ZN (N4650), .A1 (N4595), .A2 (N4531));
      NOR2_X1 XNOR_NOR2_NUM1696 (.ZN (N4654), .A1 (N4598), .A2 (N4536));
      NOR2_X1 XNOR_NOR2_NUM1697 (.ZN (N4658), .A1 (N4601), .A2 (N4541));
      NOR2_X1 XNOR_NOR2_NUM1698 (.ZN (N4662), .A1 (N4604), .A2 (N4546));
      NOR2_X1 XNOR_NOR2_NUM1699 (.ZN (N4666), .A1 (N4554), .A2 (N4607));
      NOR2_X1 XNOR_NOR2_NUM1700 (.ZN (N4667), .A1 (N4607), .A2 (N4551));
      NOR2_X1 XNOR_NOR2_NUM1701 (.ZN (N4668), .A1 (N4611), .A2 (N4612));
      NOR2_X1 XNOR_NOR2_NUM1702 (.ZN (N4671), .A1 (N4613), .A2 (N912));
      NOR2_X1 XNOR_NOR2_NUM1703 (.ZN (N4675), .A1 (N4563), .A2 (N4616));
      NOR2_X1 XNOR_NOR2_NUM1704 (.ZN (N4676), .A1 (N4616), .A2 (N960));
      NOR2_X1 XNOR_NOR2_NUM1705 (.ZN (N4677), .A1 (N4435), .A2 (N4616));
      NOR2_X1 XNOR_NOR2_NUM1706 (.ZN (N4680), .A1 (N4620), .A2 (N4621));
      NOR2_X1 XNOR_NOR2_NUM1707 (.ZN (N4683), .A1 (N4625), .A2 (N4622));
      NOR2_X1 XNOR_NOR2_NUM1708 (.ZN (N4687), .A1 (N4575), .A2 (N4628));
      NOR2_X1 XNOR_NOR2_NUM1709 (.ZN (N4688), .A1 (N4628), .A2 (N4572));
      NOR2_X1 XNOR_NOR2_NUM1710 (.ZN (N4689), .A1 (N4632), .A2 (N4633));
      NOR2_X1 XNOR_NOR2_NUM1711 (.ZN (N4692), .A1 (N4634), .A2 (N1155));
      NOR2_X1 XNOR_NOR2_NUM1712 (.ZN (N4696), .A1 (N4584), .A2 (N4637));
      NOR2_X1 XNOR_NOR2_NUM1713 (.ZN (N4697), .A1 (N4637), .A2 (N1203));
      NOR2_X1 XNOR_NOR2_NUM1714 (.ZN (N4698), .A1 (N4456), .A2 (N4637));
      NOR2_X1 XNOR_NOR2_NUM1715 (.ZN (N4701), .A1 (N4641), .A2 (N4642));
      NOR2_X1 XNOR_NOR2_NUM1716 (.ZN (N4704), .A1 (N1299), .A2 (N4643));
      NOR2_X1 XNOR_NOR2_NUM1717 (.ZN (N4708), .A1 (N4592), .A2 (N4646));
      NOR2_X1 XNOR_NOR2_NUM1718 (.ZN (N4709), .A1 (N4646), .A2 (N4526));
      NOR2_X1 XNOR_NOR2_NUM1719 (.ZN (N4710), .A1 (N4595), .A2 (N4650));
      NOR2_X1 XNOR_NOR2_NUM1720 (.ZN (N4711), .A1 (N4650), .A2 (N4531));
      NOR2_X1 XNOR_NOR2_NUM1721 (.ZN (N4712), .A1 (N4598), .A2 (N4654));
      NOR2_X1 XNOR_NOR2_NUM1722 (.ZN (N4713), .A1 (N4654), .A2 (N4536));
      NOR2_X1 XNOR_NOR2_NUM1723 (.ZN (N4714), .A1 (N4601), .A2 (N4658));
      NOR2_X1 XNOR_NOR2_NUM1724 (.ZN (N4715), .A1 (N4658), .A2 (N4541));
      NOR2_X1 XNOR_NOR2_NUM1725 (.ZN (N4716), .A1 (N4604), .A2 (N4662));
      NOR2_X1 XNOR_NOR2_NUM1726 (.ZN (N4717), .A1 (N4662), .A2 (N4546));
      NOR2_X1 XNOR_NOR2_NUM1727 (.ZN (N4718), .A1 (N4666), .A2 (N4667));
      NOR2_X1 XNOR_NOR2_NUM1728 (.ZN (N4721), .A1 (N4668), .A2 (N864));
      NOR2_X1 XNOR_NOR2_NUM1729 (.ZN (N4725), .A1 (N4613), .A2 (N4671));
      NOR2_X1 XNOR_NOR2_NUM1730 (.ZN (N4726), .A1 (N4671), .A2 (N912));
      NOR2_X1 XNOR_NOR2_NUM1731 (.ZN (N4727), .A1 (N4494), .A2 (N4671));
      NOR2_X1 XNOR_NOR2_NUM1732 (.ZN (N4730), .A1 (N4675), .A2 (N4676));
      NOR2_X1 XNOR_NOR2_NUM1733 (.ZN (N4733), .A1 (N4680), .A2 (N4677));
      NOR2_X1 XNOR_NOR2_NUM1734 (.ZN (N4737), .A1 (N4625), .A2 (N4683));
      NOR2_X1 XNOR_NOR2_NUM1735 (.ZN (N4738), .A1 (N4683), .A2 (N4622));
      NOR2_X1 XNOR_NOR2_NUM1736 (.ZN (N4739), .A1 (N4687), .A2 (N4688));
      NOR2_X1 XNOR_NOR2_NUM1737 (.ZN (N4742), .A1 (N4689), .A2 (N1107));
      NOR2_X1 XNOR_NOR2_NUM1738 (.ZN (N4746), .A1 (N4634), .A2 (N4692));
      NOR2_X1 XNOR_NOR2_NUM1739 (.ZN (N4747), .A1 (N4692), .A2 (N1155));
      NOR2_X1 XNOR_NOR2_NUM1740 (.ZN (N4748), .A1 (N4515), .A2 (N4692));
      NOR2_X1 XNOR_NOR2_NUM1741 (.ZN (N4751), .A1 (N4696), .A2 (N4697));
      NOR2_X1 XNOR_NOR2_NUM1742 (.ZN (N4754), .A1 (N4701), .A2 (N4698));
      NOR2_X1 XNOR_NOR2_NUM1743 (.ZN (N4758), .A1 (N1299), .A2 (N4704));
      NOR2_X1 XNOR_NOR2_NUM1744 (.ZN (N4759), .A1 (N4704), .A2 (N4643));
      NOR2_X1 XNOR_NOR2_NUM1745 (.ZN (N4760), .A1 (N4708), .A2 (N4709));
      NOR2_X1 XNOR_NOR2_NUM1746 (.ZN (N4763), .A1 (N4710), .A2 (N4711));
      NOR2_X1 XNOR_NOR2_NUM1747 (.ZN (N4766), .A1 (N4712), .A2 (N4713));
      NOR2_X1 XNOR_NOR2_NUM1748 (.ZN (N4769), .A1 (N4714), .A2 (N4715));
      NOR2_X1 XNOR_NOR2_NUM1749 (.ZN (N4772), .A1 (N4716), .A2 (N4717));
      NOR2_X1 XNOR_NOR2_NUM1750 (.ZN (N4775), .A1 (N4718), .A2 (N816));
      NOR2_X1 XNOR_NOR2_NUM1751 (.ZN (N4779), .A1 (N4668), .A2 (N4721));
      NOR2_X1 XNOR_NOR2_NUM1752 (.ZN (N4780), .A1 (N4721), .A2 (N864));
      NOR2_X1 XNOR_NOR2_NUM1753 (.ZN (N4781), .A1 (N4557), .A2 (N4721));
      NOR2_X1 XNOR_NOR2_NUM1754 (.ZN (N4784), .A1 (N4725), .A2 (N4726));
      NOR2_X1 XNOR_NOR2_NUM1755 (.ZN (N4787), .A1 (N4730), .A2 (N4727));
      NOR2_X1 XNOR_NOR2_NUM1756 (.ZN (N4791), .A1 (N4680), .A2 (N4733));
      NOR2_X1 XNOR_NOR2_NUM1757 (.ZN (N4792), .A1 (N4733), .A2 (N4677));
      NOR2_X1 XNOR_NOR2_NUM1758 (.ZN (N4793), .A1 (N4737), .A2 (N4738));
      NOR2_X1 XNOR_NOR2_NUM1759 (.ZN (N4796), .A1 (N4739), .A2 (N1059));
      NOR2_X1 XNOR_NOR2_NUM1760 (.ZN (N4800), .A1 (N4689), .A2 (N4742));
      NOR2_X1 XNOR_NOR2_NUM1761 (.ZN (N4801), .A1 (N4742), .A2 (N1107));
      NOR2_X1 XNOR_NOR2_NUM1762 (.ZN (N4802), .A1 (N4578), .A2 (N4742));
      NOR2_X1 XNOR_NOR2_NUM1763 (.ZN (N4805), .A1 (N4746), .A2 (N4747));
      NOR2_X1 XNOR_NOR2_NUM1764 (.ZN (N4808), .A1 (N4751), .A2 (N4748));
      NOR2_X1 XNOR_NOR2_NUM1765 (.ZN (N4812), .A1 (N4701), .A2 (N4754));
      NOR2_X1 XNOR_NOR2_NUM1766 (.ZN (N4813), .A1 (N4754), .A2 (N4698));
      NOR2_X1 XNOR_NOR2_NUM1767 (.ZN (N4814), .A1 (N4758), .A2 (N4759));
      NOR2_X1 XNOR_NOR2_NUM1768 (.ZN (N4817), .A1 (N4760), .A2 (N576));
      NOR2_X1 XNOR_NOR2_NUM1769 (.ZN (N4821), .A1 (N4763), .A2 (N624));
      NOR2_X1 XNOR_NOR2_NUM1770 (.ZN (N4825), .A1 (N4766), .A2 (N672));
      NOR2_X1 XNOR_NOR2_NUM1771 (.ZN (N4829), .A1 (N4769), .A2 (N720));
      NOR2_X1 XNOR_NOR2_NUM1772 (.ZN (N4833), .A1 (N4772), .A2 (N768));
      NOR2_X1 XNOR_NOR2_NUM1773 (.ZN (N4837), .A1 (N4718), .A2 (N4775));
      NOR2_X1 XNOR_NOR2_NUM1774 (.ZN (N4838), .A1 (N4775), .A2 (N816));
      NOR2_X1 XNOR_NOR2_NUM1775 (.ZN (N4839), .A1 (N4607), .A2 (N4775));
      NOR2_X1 XNOR_NOR2_NUM1776 (.ZN (N4842), .A1 (N4779), .A2 (N4780));
      NOR2_X1 XNOR_NOR2_NUM1777 (.ZN (N4845), .A1 (N4784), .A2 (N4781));
      NOR2_X1 XNOR_NOR2_NUM1778 (.ZN (N4849), .A1 (N4730), .A2 (N4787));
      NOR2_X1 XNOR_NOR2_NUM1779 (.ZN (N4850), .A1 (N4787), .A2 (N4727));
      NOR2_X1 XNOR_NOR2_NUM1780 (.ZN (N4851), .A1 (N4791), .A2 (N4792));
      NOR2_X1 XNOR_NOR2_NUM1781 (.ZN (N4854), .A1 (N4793), .A2 (N1011));
      NOR2_X1 XNOR_NOR2_NUM1782 (.ZN (N4858), .A1 (N4739), .A2 (N4796));
      NOR2_X1 XNOR_NOR2_NUM1783 (.ZN (N4859), .A1 (N4796), .A2 (N1059));
      NOR2_X1 XNOR_NOR2_NUM1784 (.ZN (N4860), .A1 (N4628), .A2 (N4796));
      NOR2_X1 XNOR_NOR2_NUM1785 (.ZN (N4863), .A1 (N4800), .A2 (N4801));
      NOR2_X1 XNOR_NOR2_NUM1786 (.ZN (N4866), .A1 (N4805), .A2 (N4802));
      NOR2_X1 XNOR_NOR2_NUM1787 (.ZN (N4870), .A1 (N4751), .A2 (N4808));
      NOR2_X1 XNOR_NOR2_NUM1788 (.ZN (N4871), .A1 (N4808), .A2 (N4748));
      NOR2_X1 XNOR_NOR2_NUM1789 (.ZN (N4872), .A1 (N4812), .A2 (N4813));
      NOR2_X1 XNOR_NOR2_NUM1790 (.ZN (N4875), .A1 (N4814), .A2 (N1254));
      NOR2_X1 XNOR_NOR2_NUM1791 (.ZN (N4879), .A1 (N4760), .A2 (N4817));
      NOR2_X1 XNOR_NOR2_NUM1792 (.ZN (N4880), .A1 (N4817), .A2 (N576));
      NOR2_X1 XNOR_NOR2_NUM1793 (.ZN (N4881), .A1 (N4646), .A2 (N4817));
      NOR2_X1 XNOR_NOR2_NUM1794 (.ZN (N4884), .A1 (N4763), .A2 (N4821));
      NOR2_X1 XNOR_NOR2_NUM1795 (.ZN (N4885), .A1 (N4821), .A2 (N624));
      NOR2_X1 XNOR_NOR2_NUM1796 (.ZN (N4886), .A1 (N4650), .A2 (N4821));
      NOR2_X1 XNOR_NOR2_NUM1797 (.ZN (N4889), .A1 (N4766), .A2 (N4825));
      NOR2_X1 XNOR_NOR2_NUM1798 (.ZN (N4890), .A1 (N4825), .A2 (N672));
      NOR2_X1 XNOR_NOR2_NUM1799 (.ZN (N4891), .A1 (N4654), .A2 (N4825));
      NOR2_X1 XNOR_NOR2_NUM1800 (.ZN (N4894), .A1 (N4769), .A2 (N4829));
      NOR2_X1 XNOR_NOR2_NUM1801 (.ZN (N4895), .A1 (N4829), .A2 (N720));
      NOR2_X1 XNOR_NOR2_NUM1802 (.ZN (N4896), .A1 (N4658), .A2 (N4829));
      NOR2_X1 XNOR_NOR2_NUM1803 (.ZN (N4899), .A1 (N4772), .A2 (N4833));
      NOR2_X1 XNOR_NOR2_NUM1804 (.ZN (N4900), .A1 (N4833), .A2 (N768));
      NOR2_X1 XNOR_NOR2_NUM1805 (.ZN (N4901), .A1 (N4662), .A2 (N4833));
      NOR2_X1 XNOR_NOR2_NUM1806 (.ZN (N4904), .A1 (N4837), .A2 (N4838));
      NOR2_X1 XNOR_NOR2_NUM1807 (.ZN (N4907), .A1 (N4842), .A2 (N4839));
      NOR2_X1 XNOR_NOR2_NUM1808 (.ZN (N4911), .A1 (N4784), .A2 (N4845));
      NOR2_X1 XNOR_NOR2_NUM1809 (.ZN (N4912), .A1 (N4845), .A2 (N4781));
      NOR2_X1 XNOR_NOR2_NUM1810 (.ZN (N4913), .A1 (N4849), .A2 (N4850));
      NOR2_X1 XNOR_NOR2_NUM1811 (.ZN (N4916), .A1 (N4851), .A2 (N963));
      NOR2_X1 XNOR_NOR2_NUM1812 (.ZN (N4920), .A1 (N4793), .A2 (N4854));
      NOR2_X1 XNOR_NOR2_NUM1813 (.ZN (N4921), .A1 (N4854), .A2 (N1011));
      NOR2_X1 XNOR_NOR2_NUM1814 (.ZN (N4922), .A1 (N4683), .A2 (N4854));
      NOR2_X1 XNOR_NOR2_NUM1815 (.ZN (N4925), .A1 (N4858), .A2 (N4859));
      NOR2_X1 XNOR_NOR2_NUM1816 (.ZN (N4928), .A1 (N4863), .A2 (N4860));
      NOR2_X1 XNOR_NOR2_NUM1817 (.ZN (N4932), .A1 (N4805), .A2 (N4866));
      NOR2_X1 XNOR_NOR2_NUM1818 (.ZN (N4933), .A1 (N4866), .A2 (N4802));
      NOR2_X1 XNOR_NOR2_NUM1819 (.ZN (N4934), .A1 (N4870), .A2 (N4871));
      NOR2_X1 XNOR_NOR2_NUM1820 (.ZN (N4937), .A1 (N4872), .A2 (N1206));
      NOR2_X1 XNOR_NOR2_NUM1821 (.ZN (N4941), .A1 (N4814), .A2 (N4875));
      NOR2_X1 XNOR_NOR2_NUM1822 (.ZN (N4942), .A1 (N4875), .A2 (N1254));
      NOR2_X1 XNOR_NOR2_NUM1823 (.ZN (N4943), .A1 (N4704), .A2 (N4875));
      NOR2_X1 XNOR_NOR2_NUM1824 (.ZN (N4946), .A1 (N4879), .A2 (N4880));
      NOR2_X1 XNOR_NOR2_NUM1825 (.ZN (N4947), .A1 (N4884), .A2 (N4885));
      NOR2_X1 XNOR_NOR2_NUM1826 (.ZN (N4950), .A1 (N4889), .A2 (N4890));
      NOR2_X1 XNOR_NOR2_NUM1827 (.ZN (N4953), .A1 (N4894), .A2 (N4895));
      NOR2_X1 XNOR_NOR2_NUM1828 (.ZN (N4956), .A1 (N4899), .A2 (N4900));
      NOR2_X1 XNOR_NOR2_NUM1829 (.ZN (N4959), .A1 (N4904), .A2 (N4901));
      NOR2_X1 XNOR_NOR2_NUM1830 (.ZN (N4963), .A1 (N4842), .A2 (N4907));
      NOR2_X1 XNOR_NOR2_NUM1831 (.ZN (N4964), .A1 (N4907), .A2 (N4839));
      NOR2_X1 XNOR_NOR2_NUM1832 (.ZN (N4965), .A1 (N4911), .A2 (N4912));
      NOR2_X1 XNOR_NOR2_NUM1833 (.ZN (N4968), .A1 (N4913), .A2 (N915));
      NOR2_X1 XNOR_NOR2_NUM1834 (.ZN (N4972), .A1 (N4851), .A2 (N4916));
      NOR2_X1 XNOR_NOR2_NUM1835 (.ZN (N4973), .A1 (N4916), .A2 (N963));
      NOR2_X1 XNOR_NOR2_NUM1836 (.ZN (N4974), .A1 (N4733), .A2 (N4916));
      NOR2_X1 XNOR_NOR2_NUM1837 (.ZN (N4977), .A1 (N4920), .A2 (N4921));
      NOR2_X1 XNOR_NOR2_NUM1838 (.ZN (N4980), .A1 (N4925), .A2 (N4922));
      NOR2_X1 XNOR_NOR2_NUM1839 (.ZN (N4984), .A1 (N4863), .A2 (N4928));
      NOR2_X1 XNOR_NOR2_NUM1840 (.ZN (N4985), .A1 (N4928), .A2 (N4860));
      NOR2_X1 XNOR_NOR2_NUM1841 (.ZN (N4986), .A1 (N4932), .A2 (N4933));
      NOR2_X1 XNOR_NOR2_NUM1842 (.ZN (N4989), .A1 (N4934), .A2 (N1158));
      NOR2_X1 XNOR_NOR2_NUM1843 (.ZN (N4993), .A1 (N4872), .A2 (N4937));
      NOR2_X1 XNOR_NOR2_NUM1844 (.ZN (N4994), .A1 (N4937), .A2 (N1206));
      NOR2_X1 XNOR_NOR2_NUM1845 (.ZN (N4995), .A1 (N4754), .A2 (N4937));
      NOR2_X1 XNOR_NOR2_NUM1846 (.ZN (N4998), .A1 (N4941), .A2 (N4942));
      NOR2_X1 XNOR_NOR2_NUM1847 (.ZN (N5001), .A1 (N1302), .A2 (N4943));
      NOR2_X1 XNOR_NOR2_NUM1848 (.ZN (N5005), .A1 (N4947), .A2 (N4881));
      NOR2_X1 XNOR_NOR2_NUM1849 (.ZN (N5009), .A1 (N4950), .A2 (N4886));
      NOR2_X1 XNOR_NOR2_NUM1850 (.ZN (N5013), .A1 (N4953), .A2 (N4891));
      NOR2_X1 XNOR_NOR2_NUM1851 (.ZN (N5017), .A1 (N4956), .A2 (N4896));
      NOR2_X1 XNOR_NOR2_NUM1852 (.ZN (N5021), .A1 (N4904), .A2 (N4959));
      NOR2_X1 XNOR_NOR2_NUM1853 (.ZN (N5022), .A1 (N4959), .A2 (N4901));
      NOR2_X1 XNOR_NOR2_NUM1854 (.ZN (N5023), .A1 (N4963), .A2 (N4964));
      NOR2_X1 XNOR_NOR2_NUM1855 (.ZN (N5026), .A1 (N4965), .A2 (N867));
      NOR2_X1 XNOR_NOR2_NUM1856 (.ZN (N5030), .A1 (N4913), .A2 (N4968));
      NOR2_X1 XNOR_NOR2_NUM1857 (.ZN (N5031), .A1 (N4968), .A2 (N915));
      NOR2_X1 XNOR_NOR2_NUM1858 (.ZN (N5032), .A1 (N4787), .A2 (N4968));
      NOR2_X1 XNOR_NOR2_NUM1859 (.ZN (N5035), .A1 (N4972), .A2 (N4973));
      NOR2_X1 XNOR_NOR2_NUM1860 (.ZN (N5038), .A1 (N4977), .A2 (N4974));
      NOR2_X1 XNOR_NOR2_NUM1861 (.ZN (N5042), .A1 (N4925), .A2 (N4980));
      NOR2_X1 XNOR_NOR2_NUM1862 (.ZN (N5043), .A1 (N4980), .A2 (N4922));
      NOR2_X1 XNOR_NOR2_NUM1863 (.ZN (N5044), .A1 (N4984), .A2 (N4985));
      NOR2_X1 XNOR_NOR2_NUM1864 (.ZN (N5047), .A1 (N4986), .A2 (N1110));
      NOR2_X1 XNOR_NOR2_NUM1865 (.ZN (N5051), .A1 (N4934), .A2 (N4989));
      NOR2_X1 XNOR_NOR2_NUM1866 (.ZN (N5052), .A1 (N4989), .A2 (N1158));
      NOR2_X1 XNOR_NOR2_NUM1867 (.ZN (N5053), .A1 (N4808), .A2 (N4989));
      NOR2_X1 XNOR_NOR2_NUM1868 (.ZN (N5056), .A1 (N4993), .A2 (N4994));
      NOR2_X1 XNOR_NOR2_NUM1869 (.ZN (N5059), .A1 (N4998), .A2 (N4995));
      NOR2_X1 XNOR_NOR2_NUM1870 (.ZN (N5063), .A1 (N1302), .A2 (N5001));
      NOR2_X1 XNOR_NOR2_NUM1871 (.ZN (N5064), .A1 (N5001), .A2 (N4943));
      NOR2_X1 XNOR_NOR2_NUM1872 (.ZN (N5065), .A1 (N4947), .A2 (N5005));
      NOR2_X1 XNOR_NOR2_NUM1873 (.ZN (N5066), .A1 (N5005), .A2 (N4881));
      NOR2_X1 XNOR_NOR2_NUM1874 (.ZN (N5067), .A1 (N4950), .A2 (N5009));
      NOR2_X1 XNOR_NOR2_NUM1875 (.ZN (N5068), .A1 (N5009), .A2 (N4886));
      NOR2_X1 XNOR_NOR2_NUM1876 (.ZN (N5069), .A1 (N4953), .A2 (N5013));
      NOR2_X1 XNOR_NOR2_NUM1877 (.ZN (N5070), .A1 (N5013), .A2 (N4891));
      NOR2_X1 XNOR_NOR2_NUM1878 (.ZN (N5071), .A1 (N4956), .A2 (N5017));
      NOR2_X1 XNOR_NOR2_NUM1879 (.ZN (N5072), .A1 (N5017), .A2 (N4896));
      NOR2_X1 XNOR_NOR2_NUM1880 (.ZN (N5073), .A1 (N5021), .A2 (N5022));
      NOR2_X1 XNOR_NOR2_NUM1881 (.ZN (N5076), .A1 (N5023), .A2 (N819));
      NOR2_X1 XNOR_NOR2_NUM1882 (.ZN (N5080), .A1 (N4965), .A2 (N5026));
      NOR2_X1 XNOR_NOR2_NUM1883 (.ZN (N5081), .A1 (N5026), .A2 (N867));
      NOR2_X1 XNOR_NOR2_NUM1884 (.ZN (N5082), .A1 (N4845), .A2 (N5026));
      NOR2_X1 XNOR_NOR2_NUM1885 (.ZN (N5085), .A1 (N5030), .A2 (N5031));
      NOR2_X1 XNOR_NOR2_NUM1886 (.ZN (N5088), .A1 (N5035), .A2 (N5032));
      NOR2_X1 XNOR_NOR2_NUM1887 (.ZN (N5092), .A1 (N4977), .A2 (N5038));
      NOR2_X1 XNOR_NOR2_NUM1888 (.ZN (N5093), .A1 (N5038), .A2 (N4974));
      NOR2_X1 XNOR_NOR2_NUM1889 (.ZN (N5094), .A1 (N5042), .A2 (N5043));
      NOR2_X1 XNOR_NOR2_NUM1890 (.ZN (N5097), .A1 (N5044), .A2 (N1062));
      NOR2_X1 XNOR_NOR2_NUM1891 (.ZN (N5101), .A1 (N4986), .A2 (N5047));
      NOR2_X1 XNOR_NOR2_NUM1892 (.ZN (N5102), .A1 (N5047), .A2 (N1110));
      NOR2_X1 XNOR_NOR2_NUM1893 (.ZN (N5103), .A1 (N4866), .A2 (N5047));
      NOR2_X1 XNOR_NOR2_NUM1894 (.ZN (N5106), .A1 (N5051), .A2 (N5052));
      NOR2_X1 XNOR_NOR2_NUM1895 (.ZN (N5109), .A1 (N5056), .A2 (N5053));
      NOR2_X1 XNOR_NOR2_NUM1896 (.ZN (N5113), .A1 (N4998), .A2 (N5059));
      NOR2_X1 XNOR_NOR2_NUM1897 (.ZN (N5114), .A1 (N5059), .A2 (N4995));
      NOR2_X1 XNOR_NOR2_NUM1898 (.ZN (N5115), .A1 (N5063), .A2 (N5064));
      NOR2_X1 XNOR_NOR2_NUM1899 (.ZN (N5118), .A1 (N5065), .A2 (N5066));
      NOR2_X1 XNOR_NOR2_NUM1900 (.ZN (N5121), .A1 (N5067), .A2 (N5068));
      NOR2_X1 XNOR_NOR2_NUM1901 (.ZN (N5124), .A1 (N5069), .A2 (N5070));
      NOR2_X1 XNOR_NOR2_NUM1902 (.ZN (N5127), .A1 (N5071), .A2 (N5072));
      NOR2_X1 XNOR_NOR2_NUM1903 (.ZN (N5130), .A1 (N5073), .A2 (N771));
      NOR2_X1 XNOR_NOR2_NUM1904 (.ZN (N5134), .A1 (N5023), .A2 (N5076));
      NOR2_X1 XNOR_NOR2_NUM1905 (.ZN (N5135), .A1 (N5076), .A2 (N819));
      NOR2_X1 XNOR_NOR2_NUM1906 (.ZN (N5136), .A1 (N4907), .A2 (N5076));
      NOR2_X1 XNOR_NOR2_NUM1907 (.ZN (N5139), .A1 (N5080), .A2 (N5081));
      NOR2_X1 XNOR_NOR2_NUM1908 (.ZN (N5142), .A1 (N5085), .A2 (N5082));
      NOR2_X1 XNOR_NOR2_NUM1909 (.ZN (N5146), .A1 (N5035), .A2 (N5088));
      NOR2_X1 XNOR_NOR2_NUM1910 (.ZN (N5147), .A1 (N5088), .A2 (N5032));
      NOR2_X1 XNOR_NOR2_NUM1911 (.ZN (N5148), .A1 (N5092), .A2 (N5093));
      NOR2_X1 XNOR_NOR2_NUM1912 (.ZN (N5151), .A1 (N5094), .A2 (N1014));
      NOR2_X1 XNOR_NOR2_NUM1913 (.ZN (N5155), .A1 (N5044), .A2 (N5097));
      NOR2_X1 XNOR_NOR2_NUM1914 (.ZN (N5156), .A1 (N5097), .A2 (N1062));
      NOR2_X1 XNOR_NOR2_NUM1915 (.ZN (N5157), .A1 (N4928), .A2 (N5097));
      NOR2_X1 XNOR_NOR2_NUM1916 (.ZN (N5160), .A1 (N5101), .A2 (N5102));
      NOR2_X1 XNOR_NOR2_NUM1917 (.ZN (N5163), .A1 (N5106), .A2 (N5103));
      NOR2_X1 XNOR_NOR2_NUM1918 (.ZN (N5167), .A1 (N5056), .A2 (N5109));
      NOR2_X1 XNOR_NOR2_NUM1919 (.ZN (N5168), .A1 (N5109), .A2 (N5053));
      NOR2_X1 XNOR_NOR2_NUM1920 (.ZN (N5169), .A1 (N5113), .A2 (N5114));
      NOR2_X1 XNOR_NOR2_NUM1921 (.ZN (N5172), .A1 (N5115), .A2 (N1257));
      NOR2_X1 XNOR_NOR2_NUM1922 (.ZN (N5176), .A1 (N5118), .A2 (N579));
      NOR2_X1 XNOR_NOR2_NUM1923 (.ZN (N5180), .A1 (N5121), .A2 (N627));
      NOR2_X1 XNOR_NOR2_NUM1924 (.ZN (N5184), .A1 (N5124), .A2 (N675));
      NOR2_X1 XNOR_NOR2_NUM1925 (.ZN (N5188), .A1 (N5127), .A2 (N723));
      NOR2_X1 XNOR_NOR2_NUM1926 (.ZN (N5192), .A1 (N5073), .A2 (N5130));
      NOR2_X1 XNOR_NOR2_NUM1927 (.ZN (N5193), .A1 (N5130), .A2 (N771));
      NOR2_X1 XNOR_NOR2_NUM1928 (.ZN (N5194), .A1 (N4959), .A2 (N5130));
      NOR2_X1 XNOR_NOR2_NUM1929 (.ZN (N5197), .A1 (N5134), .A2 (N5135));
      NOR2_X1 XNOR_NOR2_NUM1930 (.ZN (N5200), .A1 (N5139), .A2 (N5136));
      NOR2_X1 XNOR_NOR2_NUM1931 (.ZN (N5204), .A1 (N5085), .A2 (N5142));
      NOR2_X1 XNOR_NOR2_NUM1932 (.ZN (N5205), .A1 (N5142), .A2 (N5082));
      NOR2_X1 XNOR_NOR2_NUM1933 (.ZN (N5206), .A1 (N5146), .A2 (N5147));
      NOR2_X1 XNOR_NOR2_NUM1934 (.ZN (N5209), .A1 (N5148), .A2 (N966));
      NOR2_X1 XNOR_NOR2_NUM1935 (.ZN (N5213), .A1 (N5094), .A2 (N5151));
      NOR2_X1 XNOR_NOR2_NUM1936 (.ZN (N5214), .A1 (N5151), .A2 (N1014));
      NOR2_X1 XNOR_NOR2_NUM1937 (.ZN (N5215), .A1 (N4980), .A2 (N5151));
      NOR2_X1 XNOR_NOR2_NUM1938 (.ZN (N5218), .A1 (N5155), .A2 (N5156));
      NOR2_X1 XNOR_NOR2_NUM1939 (.ZN (N5221), .A1 (N5160), .A2 (N5157));
      NOR2_X1 XNOR_NOR2_NUM1940 (.ZN (N5225), .A1 (N5106), .A2 (N5163));
      NOR2_X1 XNOR_NOR2_NUM1941 (.ZN (N5226), .A1 (N5163), .A2 (N5103));
      NOR2_X1 XNOR_NOR2_NUM1942 (.ZN (N5227), .A1 (N5167), .A2 (N5168));
      NOR2_X1 XNOR_NOR2_NUM1943 (.ZN (N5230), .A1 (N5169), .A2 (N1209));
      NOR2_X1 XNOR_NOR2_NUM1944 (.ZN (N5234), .A1 (N5115), .A2 (N5172));
      NOR2_X1 XNOR_NOR2_NUM1945 (.ZN (N5235), .A1 (N5172), .A2 (N1257));
      NOR2_X1 XNOR_NOR2_NUM1946 (.ZN (N5236), .A1 (N5001), .A2 (N5172));
      NOR2_X1 XNOR_NOR2_NUM1947 (.ZN (N5239), .A1 (N5118), .A2 (N5176));
      NOR2_X1 XNOR_NOR2_NUM1948 (.ZN (N5240), .A1 (N5176), .A2 (N579));
      NOR2_X1 XNOR_NOR2_NUM1949 (.ZN (N5241), .A1 (N5005), .A2 (N5176));
      NOR2_X1 XNOR_NOR2_NUM1950 (.ZN (N5244), .A1 (N5121), .A2 (N5180));
      NOR2_X1 XNOR_NOR2_NUM1951 (.ZN (N5245), .A1 (N5180), .A2 (N627));
      NOR2_X1 XNOR_NOR2_NUM1952 (.ZN (N5246), .A1 (N5009), .A2 (N5180));
      NOR2_X1 XNOR_NOR2_NUM1953 (.ZN (N5249), .A1 (N5124), .A2 (N5184));
      NOR2_X1 XNOR_NOR2_NUM1954 (.ZN (N5250), .A1 (N5184), .A2 (N675));
      NOR2_X1 XNOR_NOR2_NUM1955 (.ZN (N5251), .A1 (N5013), .A2 (N5184));
      NOR2_X1 XNOR_NOR2_NUM1956 (.ZN (N5254), .A1 (N5127), .A2 (N5188));
      NOR2_X1 XNOR_NOR2_NUM1957 (.ZN (N5255), .A1 (N5188), .A2 (N723));
      NOR2_X1 XNOR_NOR2_NUM1958 (.ZN (N5256), .A1 (N5017), .A2 (N5188));
      NOR2_X1 XNOR_NOR2_NUM1959 (.ZN (N5259), .A1 (N5192), .A2 (N5193));
      NOR2_X1 XNOR_NOR2_NUM1960 (.ZN (N5262), .A1 (N5197), .A2 (N5194));
      NOR2_X1 XNOR_NOR2_NUM1961 (.ZN (N5266), .A1 (N5139), .A2 (N5200));
      NOR2_X1 XNOR_NOR2_NUM1962 (.ZN (N5267), .A1 (N5200), .A2 (N5136));
      NOR2_X1 XNOR_NOR2_NUM1963 (.ZN (N5268), .A1 (N5204), .A2 (N5205));
      NOR2_X1 XNOR_NOR2_NUM1964 (.ZN (N5271), .A1 (N5206), .A2 (N918));
      NOR2_X1 XNOR_NOR2_NUM1965 (.ZN (N5275), .A1 (N5148), .A2 (N5209));
      NOR2_X1 XNOR_NOR2_NUM1966 (.ZN (N5276), .A1 (N5209), .A2 (N966));
      NOR2_X1 XNOR_NOR2_NUM1967 (.ZN (N5277), .A1 (N5038), .A2 (N5209));
      NOR2_X1 XNOR_NOR2_NUM1968 (.ZN (N5280), .A1 (N5213), .A2 (N5214));
      NOR2_X1 XNOR_NOR2_NUM1969 (.ZN (N5283), .A1 (N5218), .A2 (N5215));
      NOR2_X1 XNOR_NOR2_NUM1970 (.ZN (N5287), .A1 (N5160), .A2 (N5221));
      NOR2_X1 XNOR_NOR2_NUM1971 (.ZN (N5288), .A1 (N5221), .A2 (N5157));
      NOR2_X1 XNOR_NOR2_NUM1972 (.ZN (N5289), .A1 (N5225), .A2 (N5226));
      NOR2_X1 XNOR_NOR2_NUM1973 (.ZN (N5292), .A1 (N5227), .A2 (N1161));
      NOR2_X1 XNOR_NOR2_NUM1974 (.ZN (N5296), .A1 (N5169), .A2 (N5230));
      NOR2_X1 XNOR_NOR2_NUM1975 (.ZN (N5297), .A1 (N5230), .A2 (N1209));
      NOR2_X1 XNOR_NOR2_NUM1976 (.ZN (N5298), .A1 (N5059), .A2 (N5230));
      NOR2_X1 XNOR_NOR2_NUM1977 (.ZN (N5301), .A1 (N5234), .A2 (N5235));
      NOR2_X1 XNOR_NOR2_NUM1978 (.ZN (N5304), .A1 (N1305), .A2 (N5236));
      NOR2_X1 XNOR_NOR2_NUM1979 (.ZN (N5308), .A1 (N5239), .A2 (N5240));
      NOR2_X1 XNOR_NOR2_NUM1980 (.ZN (N5309), .A1 (N5244), .A2 (N5245));
      NOR2_X1 XNOR_NOR2_NUM1981 (.ZN (N5312), .A1 (N5249), .A2 (N5250));
      NOR2_X1 XNOR_NOR2_NUM1982 (.ZN (N5315), .A1 (N5254), .A2 (N5255));
      NOR2_X1 XNOR_NOR2_NUM1983 (.ZN (N5318), .A1 (N5259), .A2 (N5256));
      NOR2_X1 XNOR_NOR2_NUM1984 (.ZN (N5322), .A1 (N5197), .A2 (N5262));
      NOR2_X1 XNOR_NOR2_NUM1985 (.ZN (N5323), .A1 (N5262), .A2 (N5194));
      NOR2_X1 XNOR_NOR2_NUM1986 (.ZN (N5324), .A1 (N5266), .A2 (N5267));
      NOR2_X1 XNOR_NOR2_NUM1987 (.ZN (N5327), .A1 (N5268), .A2 (N870));
      NOR2_X1 XNOR_NOR2_NUM1988 (.ZN (N5331), .A1 (N5206), .A2 (N5271));
      NOR2_X1 XNOR_NOR2_NUM1989 (.ZN (N5332), .A1 (N5271), .A2 (N918));
      NOR2_X1 XNOR_NOR2_NUM1990 (.ZN (N5333), .A1 (N5088), .A2 (N5271));
      NOR2_X1 XNOR_NOR2_NUM1991 (.ZN (N5336), .A1 (N5275), .A2 (N5276));
      NOR2_X1 XNOR_NOR2_NUM1992 (.ZN (N5339), .A1 (N5280), .A2 (N5277));
      NOR2_X1 XNOR_NOR2_NUM1993 (.ZN (N5343), .A1 (N5218), .A2 (N5283));
      NOR2_X1 XNOR_NOR2_NUM1994 (.ZN (N5344), .A1 (N5283), .A2 (N5215));
      NOR2_X1 XNOR_NOR2_NUM1995 (.ZN (N5345), .A1 (N5287), .A2 (N5288));
      NOR2_X1 XNOR_NOR2_NUM1996 (.ZN (N5348), .A1 (N5289), .A2 (N1113));
      NOR2_X1 XNOR_NOR2_NUM1997 (.ZN (N5352), .A1 (N5227), .A2 (N5292));
      NOR2_X1 XNOR_NOR2_NUM1998 (.ZN (N5353), .A1 (N5292), .A2 (N1161));
      NOR2_X1 XNOR_NOR2_NUM1999 (.ZN (N5354), .A1 (N5109), .A2 (N5292));
      NOR2_X1 XNOR_NOR2_NUM2000 (.ZN (N5357), .A1 (N5296), .A2 (N5297));
      NOR2_X1 XNOR_NOR2_NUM2001 (.ZN (N5360), .A1 (N5301), .A2 (N5298));
      NOR2_X1 XNOR_NOR2_NUM2002 (.ZN (N5364), .A1 (N1305), .A2 (N5304));
      NOR2_X1 XNOR_NOR2_NUM2003 (.ZN (N5365), .A1 (N5304), .A2 (N5236));
      NOR2_X1 XNOR_NOR2_NUM2004 (.ZN (N5366), .A1 (N5309), .A2 (N5241));
      NOR2_X1 XNOR_NOR2_NUM2005 (.ZN (N5370), .A1 (N5312), .A2 (N5246));
      NOR2_X1 XNOR_NOR2_NUM2006 (.ZN (N5374), .A1 (N5315), .A2 (N5251));
      NOR2_X1 XNOR_NOR2_NUM2007 (.ZN (N5378), .A1 (N5259), .A2 (N5318));
      NOR2_X1 XNOR_NOR2_NUM2008 (.ZN (N5379), .A1 (N5318), .A2 (N5256));
      NOR2_X1 XNOR_NOR2_NUM2009 (.ZN (N5380), .A1 (N5322), .A2 (N5323));
      NOR2_X1 XNOR_NOR2_NUM2010 (.ZN (N5383), .A1 (N5324), .A2 (N822));
      NOR2_X1 XNOR_NOR2_NUM2011 (.ZN (N5387), .A1 (N5268), .A2 (N5327));
      NOR2_X1 XNOR_NOR2_NUM2012 (.ZN (N5388), .A1 (N5327), .A2 (N870));
      NOR2_X1 XNOR_NOR2_NUM2013 (.ZN (N5389), .A1 (N5142), .A2 (N5327));
      NOR2_X1 XNOR_NOR2_NUM2014 (.ZN (N5392), .A1 (N5331), .A2 (N5332));
      NOR2_X1 XNOR_NOR2_NUM2015 (.ZN (N5395), .A1 (N5336), .A2 (N5333));
      NOR2_X1 XNOR_NOR2_NUM2016 (.ZN (N5399), .A1 (N5280), .A2 (N5339));
      NOR2_X1 XNOR_NOR2_NUM2017 (.ZN (N5400), .A1 (N5339), .A2 (N5277));
      NOR2_X1 XNOR_NOR2_NUM2018 (.ZN (N5401), .A1 (N5343), .A2 (N5344));
      NOR2_X1 XNOR_NOR2_NUM2019 (.ZN (N5404), .A1 (N5345), .A2 (N1065));
      NOR2_X1 XNOR_NOR2_NUM2020 (.ZN (N5408), .A1 (N5289), .A2 (N5348));
      NOR2_X1 XNOR_NOR2_NUM2021 (.ZN (N5409), .A1 (N5348), .A2 (N1113));
      NOR2_X1 XNOR_NOR2_NUM2022 (.ZN (N5410), .A1 (N5163), .A2 (N5348));
      NOR2_X1 XNOR_NOR2_NUM2023 (.ZN (N5413), .A1 (N5352), .A2 (N5353));
      NOR2_X1 XNOR_NOR2_NUM2024 (.ZN (N5416), .A1 (N5357), .A2 (N5354));
      NOR2_X1 XNOR_NOR2_NUM2025 (.ZN (N5420), .A1 (N5301), .A2 (N5360));
      NOR2_X1 XNOR_NOR2_NUM2026 (.ZN (N5421), .A1 (N5360), .A2 (N5298));
      NOR2_X1 XNOR_NOR2_NUM2027 (.ZN (N5422), .A1 (N5364), .A2 (N5365));
      NOR2_X1 XNOR_NOR2_NUM2028 (.ZN (N5425), .A1 (N5309), .A2 (N5366));
      NOR2_X1 XNOR_NOR2_NUM2029 (.ZN (N5426), .A1 (N5366), .A2 (N5241));
      NOR2_X1 XNOR_NOR2_NUM2030 (.ZN (N5427), .A1 (N5312), .A2 (N5370));
      NOR2_X1 XNOR_NOR2_NUM2031 (.ZN (N5428), .A1 (N5370), .A2 (N5246));
      NOR2_X1 XNOR_NOR2_NUM2032 (.ZN (N5429), .A1 (N5315), .A2 (N5374));
      NOR2_X1 XNOR_NOR2_NUM2033 (.ZN (N5430), .A1 (N5374), .A2 (N5251));
      NOR2_X1 XNOR_NOR2_NUM2034 (.ZN (N5431), .A1 (N5378), .A2 (N5379));
      NOR2_X1 XNOR_NOR2_NUM2035 (.ZN (N5434), .A1 (N5380), .A2 (N774));
      NOR2_X1 XNOR_NOR2_NUM2036 (.ZN (N5438), .A1 (N5324), .A2 (N5383));
      NOR2_X1 XNOR_NOR2_NUM2037 (.ZN (N5439), .A1 (N5383), .A2 (N822));
      NOR2_X1 XNOR_NOR2_NUM2038 (.ZN (N5440), .A1 (N5200), .A2 (N5383));
      NOR2_X1 XNOR_NOR2_NUM2039 (.ZN (N5443), .A1 (N5387), .A2 (N5388));
      NOR2_X1 XNOR_NOR2_NUM2040 (.ZN (N5446), .A1 (N5392), .A2 (N5389));
      NOR2_X1 XNOR_NOR2_NUM2041 (.ZN (N5450), .A1 (N5336), .A2 (N5395));
      NOR2_X1 XNOR_NOR2_NUM2042 (.ZN (N5451), .A1 (N5395), .A2 (N5333));
      NOR2_X1 XNOR_NOR2_NUM2043 (.ZN (N5452), .A1 (N5399), .A2 (N5400));
      NOR2_X1 XNOR_NOR2_NUM2044 (.ZN (N5455), .A1 (N5401), .A2 (N1017));
      NOR2_X1 XNOR_NOR2_NUM2045 (.ZN (N5459), .A1 (N5345), .A2 (N5404));
      NOR2_X1 XNOR_NOR2_NUM2046 (.ZN (N5460), .A1 (N5404), .A2 (N1065));
      NOR2_X1 XNOR_NOR2_NUM2047 (.ZN (N5461), .A1 (N5221), .A2 (N5404));
      NOR2_X1 XNOR_NOR2_NUM2048 (.ZN (N5464), .A1 (N5408), .A2 (N5409));
      NOR2_X1 XNOR_NOR2_NUM2049 (.ZN (N5467), .A1 (N5413), .A2 (N5410));
      NOR2_X1 XNOR_NOR2_NUM2050 (.ZN (N5471), .A1 (N5357), .A2 (N5416));
      NOR2_X1 XNOR_NOR2_NUM2051 (.ZN (N5472), .A1 (N5416), .A2 (N5354));
      NOR2_X1 XNOR_NOR2_NUM2052 (.ZN (N5473), .A1 (N5420), .A2 (N5421));
      NOR2_X1 XNOR_NOR2_NUM2053 (.ZN (N5476), .A1 (N5422), .A2 (N1260));
      NOR2_X1 XNOR_NOR2_NUM2054 (.ZN (N5480), .A1 (N5425), .A2 (N5426));
      NOR2_X1 XNOR_NOR2_NUM2055 (.ZN (N5483), .A1 (N5427), .A2 (N5428));
      NOR2_X1 XNOR_NOR2_NUM2056 (.ZN (N5486), .A1 (N5429), .A2 (N5430));
      NOR2_X1 XNOR_NOR2_NUM2057 (.ZN (N5489), .A1 (N5431), .A2 (N726));
      NOR2_X1 XNOR_NOR2_NUM2058 (.ZN (N5493), .A1 (N5380), .A2 (N5434));
      NOR2_X1 XNOR_NOR2_NUM2059 (.ZN (N5494), .A1 (N5434), .A2 (N774));
      NOR2_X1 XNOR_NOR2_NUM2060 (.ZN (N5495), .A1 (N5262), .A2 (N5434));
      NOR2_X1 XNOR_NOR2_NUM2061 (.ZN (N5498), .A1 (N5438), .A2 (N5439));
      NOR2_X1 XNOR_NOR2_NUM2062 (.ZN (N5501), .A1 (N5443), .A2 (N5440));
      NOR2_X1 XNOR_NOR2_NUM2063 (.ZN (N5505), .A1 (N5392), .A2 (N5446));
      NOR2_X1 XNOR_NOR2_NUM2064 (.ZN (N5506), .A1 (N5446), .A2 (N5389));
      NOR2_X1 XNOR_NOR2_NUM2065 (.ZN (N5507), .A1 (N5450), .A2 (N5451));
      NOR2_X1 XNOR_NOR2_NUM2066 (.ZN (N5510), .A1 (N5452), .A2 (N969));
      NOR2_X1 XNOR_NOR2_NUM2067 (.ZN (N5514), .A1 (N5401), .A2 (N5455));
      NOR2_X1 XNOR_NOR2_NUM2068 (.ZN (N5515), .A1 (N5455), .A2 (N1017));
      NOR2_X1 XNOR_NOR2_NUM2069 (.ZN (N5516), .A1 (N5283), .A2 (N5455));
      NOR2_X1 XNOR_NOR2_NUM2070 (.ZN (N5519), .A1 (N5459), .A2 (N5460));
      NOR2_X1 XNOR_NOR2_NUM2071 (.ZN (N5522), .A1 (N5464), .A2 (N5461));
      NOR2_X1 XNOR_NOR2_NUM2072 (.ZN (N5526), .A1 (N5413), .A2 (N5467));
      NOR2_X1 XNOR_NOR2_NUM2073 (.ZN (N5527), .A1 (N5467), .A2 (N5410));
      NOR2_X1 XNOR_NOR2_NUM2074 (.ZN (N5528), .A1 (N5471), .A2 (N5472));
      NOR2_X1 XNOR_NOR2_NUM2075 (.ZN (N5531), .A1 (N5473), .A2 (N1212));
      NOR2_X1 XNOR_NOR2_NUM2076 (.ZN (N5535), .A1 (N5422), .A2 (N5476));
      NOR2_X1 XNOR_NOR2_NUM2077 (.ZN (N5536), .A1 (N5476), .A2 (N1260));
      NOR2_X1 XNOR_NOR2_NUM2078 (.ZN (N5537), .A1 (N5304), .A2 (N5476));
      NOR2_X1 XNOR_NOR2_NUM2079 (.ZN (N5540), .A1 (N5480), .A2 (N582));
      NOR2_X1 XNOR_NOR2_NUM2080 (.ZN (N5544), .A1 (N5483), .A2 (N630));
      NOR2_X1 XNOR_NOR2_NUM2081 (.ZN (N5548), .A1 (N5486), .A2 (N678));
      NOR2_X1 XNOR_NOR2_NUM2082 (.ZN (N5552), .A1 (N5431), .A2 (N5489));
      NOR2_X1 XNOR_NOR2_NUM2083 (.ZN (N5553), .A1 (N5489), .A2 (N726));
      NOR2_X1 XNOR_NOR2_NUM2084 (.ZN (N5554), .A1 (N5318), .A2 (N5489));
      NOR2_X1 XNOR_NOR2_NUM2085 (.ZN (N5557), .A1 (N5493), .A2 (N5494));
      NOR2_X1 XNOR_NOR2_NUM2086 (.ZN (N5560), .A1 (N5498), .A2 (N5495));
      NOR2_X1 XNOR_NOR2_NUM2087 (.ZN (N5564), .A1 (N5443), .A2 (N5501));
      NOR2_X1 XNOR_NOR2_NUM2088 (.ZN (N5565), .A1 (N5501), .A2 (N5440));
      NOR2_X1 XNOR_NOR2_NUM2089 (.ZN (N5566), .A1 (N5505), .A2 (N5506));
      NOR2_X1 XNOR_NOR2_NUM2090 (.ZN (N5569), .A1 (N5507), .A2 (N921));
      NOR2_X1 XNOR_NOR2_NUM2091 (.ZN (N5573), .A1 (N5452), .A2 (N5510));
      NOR2_X1 XNOR_NOR2_NUM2092 (.ZN (N5574), .A1 (N5510), .A2 (N969));
      NOR2_X1 XNOR_NOR2_NUM2093 (.ZN (N5575), .A1 (N5339), .A2 (N5510));
      NOR2_X1 XNOR_NOR2_NUM2094 (.ZN (N5578), .A1 (N5514), .A2 (N5515));
      NOR2_X1 XNOR_NOR2_NUM2095 (.ZN (N5581), .A1 (N5519), .A2 (N5516));
      NOR2_X1 XNOR_NOR2_NUM2096 (.ZN (N5585), .A1 (N5464), .A2 (N5522));
      NOR2_X1 XNOR_NOR2_NUM2097 (.ZN (N5586), .A1 (N5522), .A2 (N5461));
      NOR2_X1 XNOR_NOR2_NUM2098 (.ZN (N5587), .A1 (N5526), .A2 (N5527));
      NOR2_X1 XNOR_NOR2_NUM2099 (.ZN (N5590), .A1 (N5528), .A2 (N1164));
      NOR2_X1 XNOR_NOR2_NUM2100 (.ZN (N5594), .A1 (N5473), .A2 (N5531));
      NOR2_X1 XNOR_NOR2_NUM2101 (.ZN (N5595), .A1 (N5531), .A2 (N1212));
      NOR2_X1 XNOR_NOR2_NUM2102 (.ZN (N5596), .A1 (N5360), .A2 (N5531));
      NOR2_X1 XNOR_NOR2_NUM2103 (.ZN (N5599), .A1 (N5535), .A2 (N5536));
      NOR2_X1 XNOR_NOR2_NUM2104 (.ZN (N5602), .A1 (N1308), .A2 (N5537));
      NOR2_X1 XNOR_NOR2_NUM2105 (.ZN (N5606), .A1 (N5480), .A2 (N5540));
      NOR2_X1 XNOR_NOR2_NUM2106 (.ZN (N5607), .A1 (N5540), .A2 (N582));
      NOR2_X1 XNOR_NOR2_NUM2107 (.ZN (N5608), .A1 (N5366), .A2 (N5540));
      NOR2_X1 XNOR_NOR2_NUM2108 (.ZN (N5611), .A1 (N5483), .A2 (N5544));
      NOR2_X1 XNOR_NOR2_NUM2109 (.ZN (N5612), .A1 (N5544), .A2 (N630));
      NOR2_X1 XNOR_NOR2_NUM2110 (.ZN (N5613), .A1 (N5370), .A2 (N5544));
      NOR2_X1 XNOR_NOR2_NUM2111 (.ZN (N5616), .A1 (N5486), .A2 (N5548));
      NOR2_X1 XNOR_NOR2_NUM2112 (.ZN (N5617), .A1 (N5548), .A2 (N678));
      NOR2_X1 XNOR_NOR2_NUM2113 (.ZN (N5618), .A1 (N5374), .A2 (N5548));
      NOR2_X1 XNOR_NOR2_NUM2114 (.ZN (N5621), .A1 (N5552), .A2 (N5553));
      NOR2_X1 XNOR_NOR2_NUM2115 (.ZN (N5624), .A1 (N5557), .A2 (N5554));
      NOR2_X1 XNOR_NOR2_NUM2116 (.ZN (N5628), .A1 (N5498), .A2 (N5560));
      NOR2_X1 XNOR_NOR2_NUM2117 (.ZN (N5629), .A1 (N5560), .A2 (N5495));
      NOR2_X1 XNOR_NOR2_NUM2118 (.ZN (N5630), .A1 (N5564), .A2 (N5565));
      NOR2_X1 XNOR_NOR2_NUM2119 (.ZN (N5633), .A1 (N5566), .A2 (N873));
      NOR2_X1 XNOR_NOR2_NUM2120 (.ZN (N5637), .A1 (N5507), .A2 (N5569));
      NOR2_X1 XNOR_NOR2_NUM2121 (.ZN (N5638), .A1 (N5569), .A2 (N921));
      NOR2_X1 XNOR_NOR2_NUM2122 (.ZN (N5639), .A1 (N5395), .A2 (N5569));
      NOR2_X1 XNOR_NOR2_NUM2123 (.ZN (N5642), .A1 (N5573), .A2 (N5574));
      NOR2_X1 XNOR_NOR2_NUM2124 (.ZN (N5645), .A1 (N5578), .A2 (N5575));
      NOR2_X1 XNOR_NOR2_NUM2125 (.ZN (N5649), .A1 (N5519), .A2 (N5581));
      NOR2_X1 XNOR_NOR2_NUM2126 (.ZN (N5650), .A1 (N5581), .A2 (N5516));
      NOR2_X1 XNOR_NOR2_NUM2127 (.ZN (N5651), .A1 (N5585), .A2 (N5586));
      NOR2_X1 XNOR_NOR2_NUM2128 (.ZN (N5654), .A1 (N5587), .A2 (N1116));
      NOR2_X1 XNOR_NOR2_NUM2129 (.ZN (N5658), .A1 (N5528), .A2 (N5590));
      NOR2_X1 XNOR_NOR2_NUM2130 (.ZN (N5659), .A1 (N5590), .A2 (N1164));
      NOR2_X1 XNOR_NOR2_NUM2131 (.ZN (N5660), .A1 (N5416), .A2 (N5590));
      NOR2_X1 XNOR_NOR2_NUM2132 (.ZN (N5663), .A1 (N5594), .A2 (N5595));
      NOR2_X1 XNOR_NOR2_NUM2133 (.ZN (N5666), .A1 (N5599), .A2 (N5596));
      NOR2_X1 XNOR_NOR2_NUM2134 (.ZN (N5670), .A1 (N1308), .A2 (N5602));
      NOR2_X1 XNOR_NOR2_NUM2135 (.ZN (N5671), .A1 (N5602), .A2 (N5537));
      NOR2_X1 XNOR_NOR2_NUM2136 (.ZN (N5672), .A1 (N5606), .A2 (N5607));
      NOR2_X1 XNOR_NOR2_NUM2137 (.ZN (N5673), .A1 (N5611), .A2 (N5612));
      NOR2_X1 XNOR_NOR2_NUM2138 (.ZN (N5676), .A1 (N5616), .A2 (N5617));
      NOR2_X1 XNOR_NOR2_NUM2139 (.ZN (N5679), .A1 (N5621), .A2 (N5618));
      NOR2_X1 XNOR_NOR2_NUM2140 (.ZN (N5683), .A1 (N5557), .A2 (N5624));
      NOR2_X1 XNOR_NOR2_NUM2141 (.ZN (N5684), .A1 (N5624), .A2 (N5554));
      NOR2_X1 XNOR_NOR2_NUM2142 (.ZN (N5685), .A1 (N5628), .A2 (N5629));
      NOR2_X1 XNOR_NOR2_NUM2143 (.ZN (N5688), .A1 (N5630), .A2 (N825));
      NOR2_X1 XNOR_NOR2_NUM2144 (.ZN (N5692), .A1 (N5566), .A2 (N5633));
      NOR2_X1 XNOR_NOR2_NUM2145 (.ZN (N5693), .A1 (N5633), .A2 (N873));
      NOR2_X1 XNOR_NOR2_NUM2146 (.ZN (N5694), .A1 (N5446), .A2 (N5633));
      NOR2_X1 XNOR_NOR2_NUM2147 (.ZN (N5697), .A1 (N5637), .A2 (N5638));
      NOR2_X1 XNOR_NOR2_NUM2148 (.ZN (N5700), .A1 (N5642), .A2 (N5639));
      NOR2_X1 XNOR_NOR2_NUM2149 (.ZN (N5704), .A1 (N5578), .A2 (N5645));
      NOR2_X1 XNOR_NOR2_NUM2150 (.ZN (N5705), .A1 (N5645), .A2 (N5575));
      NOR2_X1 XNOR_NOR2_NUM2151 (.ZN (N5706), .A1 (N5649), .A2 (N5650));
      NOR2_X1 XNOR_NOR2_NUM2152 (.ZN (N5709), .A1 (N5651), .A2 (N1068));
      NOR2_X1 XNOR_NOR2_NUM2153 (.ZN (N5713), .A1 (N5587), .A2 (N5654));
      NOR2_X1 XNOR_NOR2_NUM2154 (.ZN (N5714), .A1 (N5654), .A2 (N1116));
      NOR2_X1 XNOR_NOR2_NUM2155 (.ZN (N5715), .A1 (N5467), .A2 (N5654));
      NOR2_X1 XNOR_NOR2_NUM2156 (.ZN (N5718), .A1 (N5658), .A2 (N5659));
      NOR2_X1 XNOR_NOR2_NUM2157 (.ZN (N5721), .A1 (N5663), .A2 (N5660));
      NOR2_X1 XNOR_NOR2_NUM2158 (.ZN (N5725), .A1 (N5599), .A2 (N5666));
      NOR2_X1 XNOR_NOR2_NUM2159 (.ZN (N5726), .A1 (N5666), .A2 (N5596));
      NOR2_X1 XNOR_NOR2_NUM2160 (.ZN (N5727), .A1 (N5670), .A2 (N5671));
      NOR2_X1 XNOR_NOR2_NUM2161 (.ZN (N5730), .A1 (N5673), .A2 (N5608));
      NOR2_X1 XNOR_NOR2_NUM2162 (.ZN (N5734), .A1 (N5676), .A2 (N5613));
      NOR2_X1 XNOR_NOR2_NUM2163 (.ZN (N5738), .A1 (N5621), .A2 (N5679));
      NOR2_X1 XNOR_NOR2_NUM2164 (.ZN (N5739), .A1 (N5679), .A2 (N5618));
      NOR2_X1 XNOR_NOR2_NUM2165 (.ZN (N5740), .A1 (N5683), .A2 (N5684));
      NOR2_X1 XNOR_NOR2_NUM2166 (.ZN (N5743), .A1 (N5685), .A2 (N777));
      NOR2_X1 XNOR_NOR2_NUM2167 (.ZN (N5747), .A1 (N5630), .A2 (N5688));
      NOR2_X1 XNOR_NOR2_NUM2168 (.ZN (N5748), .A1 (N5688), .A2 (N825));
      NOR2_X1 XNOR_NOR2_NUM2169 (.ZN (N5749), .A1 (N5501), .A2 (N5688));
      NOR2_X1 XNOR_NOR2_NUM2170 (.ZN (N5752), .A1 (N5692), .A2 (N5693));
      NOR2_X1 XNOR_NOR2_NUM2171 (.ZN (N5755), .A1 (N5697), .A2 (N5694));
      NOR2_X1 XNOR_NOR2_NUM2172 (.ZN (N5759), .A1 (N5642), .A2 (N5700));
      NOR2_X1 XNOR_NOR2_NUM2173 (.ZN (N5760), .A1 (N5700), .A2 (N5639));
      NOR2_X1 XNOR_NOR2_NUM2174 (.ZN (N5761), .A1 (N5704), .A2 (N5705));
      NOR2_X1 XNOR_NOR2_NUM2175 (.ZN (N5764), .A1 (N5706), .A2 (N1020));
      NOR2_X1 XNOR_NOR2_NUM2176 (.ZN (N5768), .A1 (N5651), .A2 (N5709));
      NOR2_X1 XNOR_NOR2_NUM2177 (.ZN (N5769), .A1 (N5709), .A2 (N1068));
      NOR2_X1 XNOR_NOR2_NUM2178 (.ZN (N5770), .A1 (N5522), .A2 (N5709));
      NOR2_X1 XNOR_NOR2_NUM2179 (.ZN (N5773), .A1 (N5713), .A2 (N5714));
      NOR2_X1 XNOR_NOR2_NUM2180 (.ZN (N5776), .A1 (N5718), .A2 (N5715));
      NOR2_X1 XNOR_NOR2_NUM2181 (.ZN (N5780), .A1 (N5663), .A2 (N5721));
      NOR2_X1 XNOR_NOR2_NUM2182 (.ZN (N5781), .A1 (N5721), .A2 (N5660));
      NOR2_X1 XNOR_NOR2_NUM2183 (.ZN (N5782), .A1 (N5725), .A2 (N5726));
      NOR2_X1 XNOR_NOR2_NUM2184 (.ZN (N5785), .A1 (N5673), .A2 (N5730));
      NOR2_X1 XNOR_NOR2_NUM2185 (.ZN (N5786), .A1 (N5730), .A2 (N5608));
      NOR2_X1 XNOR_NOR2_NUM2186 (.ZN (N5787), .A1 (N5676), .A2 (N5734));
      NOR2_X1 XNOR_NOR2_NUM2187 (.ZN (N5788), .A1 (N5734), .A2 (N5613));
      NOR2_X1 XNOR_NOR2_NUM2188 (.ZN (N5789), .A1 (N5738), .A2 (N5739));
      NOR2_X1 XNOR_NOR2_NUM2189 (.ZN (N5792), .A1 (N5740), .A2 (N729));
      NOR2_X1 XNOR_NOR2_NUM2190 (.ZN (N5796), .A1 (N5685), .A2 (N5743));
      NOR2_X1 XNOR_NOR2_NUM2191 (.ZN (N5797), .A1 (N5743), .A2 (N777));
      NOR2_X1 XNOR_NOR2_NUM2192 (.ZN (N5798), .A1 (N5560), .A2 (N5743));
      NOR2_X1 XNOR_NOR2_NUM2193 (.ZN (N5801), .A1 (N5747), .A2 (N5748));
      NOR2_X1 XNOR_NOR2_NUM2194 (.ZN (N5804), .A1 (N5752), .A2 (N5749));
      NOR2_X1 XNOR_NOR2_NUM2195 (.ZN (N5808), .A1 (N5697), .A2 (N5755));
      NOR2_X1 XNOR_NOR2_NUM2196 (.ZN (N5809), .A1 (N5755), .A2 (N5694));
      NOR2_X1 XNOR_NOR2_NUM2197 (.ZN (N5810), .A1 (N5759), .A2 (N5760));
      NOR2_X1 XNOR_NOR2_NUM2198 (.ZN (N5813), .A1 (N5761), .A2 (N972));
      NOR2_X1 XNOR_NOR2_NUM2199 (.ZN (N5817), .A1 (N5706), .A2 (N5764));
      NOR2_X1 XNOR_NOR2_NUM2200 (.ZN (N5818), .A1 (N5764), .A2 (N1020));
      NOR2_X1 XNOR_NOR2_NUM2201 (.ZN (N5819), .A1 (N5581), .A2 (N5764));
      NOR2_X1 XNOR_NOR2_NUM2202 (.ZN (N5822), .A1 (N5768), .A2 (N5769));
      NOR2_X1 XNOR_NOR2_NUM2203 (.ZN (N5825), .A1 (N5773), .A2 (N5770));
      NOR2_X1 XNOR_NOR2_NUM2204 (.ZN (N5829), .A1 (N5718), .A2 (N5776));
      NOR2_X1 XNOR_NOR2_NUM2205 (.ZN (N5830), .A1 (N5776), .A2 (N5715));
      NOR2_X1 XNOR_NOR2_NUM2206 (.ZN (N5831), .A1 (N5780), .A2 (N5781));
      NOR2_X1 XNOR_NOR2_NUM2207 (.ZN (N5834), .A1 (N5785), .A2 (N5786));
      NOR2_X1 XNOR_NOR2_NUM2208 (.ZN (N5837), .A1 (N5787), .A2 (N5788));
      NOR2_X1 XNOR_NOR2_NUM2209 (.ZN (N5840), .A1 (N5789), .A2 (N681));
      NOR2_X1 XNOR_NOR2_NUM2210 (.ZN (N5844), .A1 (N5740), .A2 (N5792));
      NOR2_X1 XNOR_NOR2_NUM2211 (.ZN (N5845), .A1 (N5792), .A2 (N729));
      NOR2_X1 XNOR_NOR2_NUM2212 (.ZN (N5846), .A1 (N5624), .A2 (N5792));
      NOR2_X1 XNOR_NOR2_NUM2213 (.ZN (N5849), .A1 (N5796), .A2 (N5797));
      NOR2_X1 XNOR_NOR2_NUM2214 (.ZN (N5852), .A1 (N5801), .A2 (N5798));
      NOR2_X1 XNOR_NOR2_NUM2215 (.ZN (N5856), .A1 (N5752), .A2 (N5804));
      NOR2_X1 XNOR_NOR2_NUM2216 (.ZN (N5857), .A1 (N5804), .A2 (N5749));
      NOR2_X1 XNOR_NOR2_NUM2217 (.ZN (N5858), .A1 (N5808), .A2 (N5809));
      NOR2_X1 XNOR_NOR2_NUM2218 (.ZN (N5861), .A1 (N5810), .A2 (N924));
      NOR2_X1 XNOR_NOR2_NUM2219 (.ZN (N5865), .A1 (N5761), .A2 (N5813));
      NOR2_X1 XNOR_NOR2_NUM2220 (.ZN (N5866), .A1 (N5813), .A2 (N972));
      NOR2_X1 XNOR_NOR2_NUM2221 (.ZN (N5867), .A1 (N5645), .A2 (N5813));
      NOR2_X1 XNOR_NOR2_NUM2222 (.ZN (N5870), .A1 (N5817), .A2 (N5818));
      NOR2_X1 XNOR_NOR2_NUM2223 (.ZN (N5873), .A1 (N5822), .A2 (N5819));
      NOR2_X1 XNOR_NOR2_NUM2224 (.ZN (N5877), .A1 (N5773), .A2 (N5825));
      NOR2_X1 XNOR_NOR2_NUM2225 (.ZN (N5878), .A1 (N5825), .A2 (N5770));
      NOR2_X1 XNOR_NOR2_NUM2226 (.ZN (N5879), .A1 (N5829), .A2 (N5830));
      NOR2_X1 XNOR_NOR2_NUM2227 (.ZN (N5882), .A1 (N5834), .A2 (N585));
      NOR2_X1 XNOR_NOR2_NUM2228 (.ZN (N5886), .A1 (N5837), .A2 (N633));
      NOR2_X1 XNOR_NOR2_NUM2229 (.ZN (N5890), .A1 (N5789), .A2 (N5840));
      NOR2_X1 XNOR_NOR2_NUM2230 (.ZN (N5891), .A1 (N5840), .A2 (N681));
      NOR2_X1 XNOR_NOR2_NUM2231 (.ZN (N5892), .A1 (N5679), .A2 (N5840));
      NOR2_X1 XNOR_NOR2_NUM2232 (.ZN (N5895), .A1 (N5844), .A2 (N5845));
      NOR2_X1 XNOR_NOR2_NUM2233 (.ZN (N5898), .A1 (N5849), .A2 (N5846));
      NOR2_X1 XNOR_NOR2_NUM2234 (.ZN (N5902), .A1 (N5801), .A2 (N5852));
      NOR2_X1 XNOR_NOR2_NUM2235 (.ZN (N5903), .A1 (N5852), .A2 (N5798));
      NOR2_X1 XNOR_NOR2_NUM2236 (.ZN (N5904), .A1 (N5856), .A2 (N5857));
      NOR2_X1 XNOR_NOR2_NUM2237 (.ZN (N5907), .A1 (N5858), .A2 (N876));
      NOR2_X1 XNOR_NOR2_NUM2238 (.ZN (N5911), .A1 (N5810), .A2 (N5861));
      NOR2_X1 XNOR_NOR2_NUM2239 (.ZN (N5912), .A1 (N5861), .A2 (N924));
      NOR2_X1 XNOR_NOR2_NUM2240 (.ZN (N5913), .A1 (N5700), .A2 (N5861));
      NOR2_X1 XNOR_NOR2_NUM2241 (.ZN (N5916), .A1 (N5865), .A2 (N5866));
      NOR2_X1 XNOR_NOR2_NUM2242 (.ZN (N5919), .A1 (N5870), .A2 (N5867));
      NOR2_X1 XNOR_NOR2_NUM2243 (.ZN (N5923), .A1 (N5822), .A2 (N5873));
      NOR2_X1 XNOR_NOR2_NUM2244 (.ZN (N5924), .A1 (N5873), .A2 (N5819));
      NOR2_X1 XNOR_NOR2_NUM2245 (.ZN (N5925), .A1 (N5877), .A2 (N5878));
      NOR2_X1 XNOR_NOR2_NUM2246 (.ZN (N5928), .A1 (N5834), .A2 (N5882));
      NOR2_X1 XNOR_NOR2_NUM2247 (.ZN (N5929), .A1 (N5882), .A2 (N585));
      NOR2_X1 XNOR_NOR2_NUM2248 (.ZN (N5930), .A1 (N5730), .A2 (N5882));
      NOR2_X1 XNOR_NOR2_NUM2249 (.ZN (N5933), .A1 (N5837), .A2 (N5886));
      NOR2_X1 XNOR_NOR2_NUM2250 (.ZN (N5934), .A1 (N5886), .A2 (N633));
      NOR2_X1 XNOR_NOR2_NUM2251 (.ZN (N5935), .A1 (N5734), .A2 (N5886));
      NOR2_X1 XNOR_NOR2_NUM2252 (.ZN (N5938), .A1 (N5890), .A2 (N5891));
      NOR2_X1 XNOR_NOR2_NUM2253 (.ZN (N5941), .A1 (N5895), .A2 (N5892));
      NOR2_X1 XNOR_NOR2_NUM2254 (.ZN (N5945), .A1 (N5849), .A2 (N5898));
      NOR2_X1 XNOR_NOR2_NUM2255 (.ZN (N5946), .A1 (N5898), .A2 (N5846));
      NOR2_X1 XNOR_NOR2_NUM2256 (.ZN (N5947), .A1 (N5902), .A2 (N5903));
      NOR2_X1 XNOR_NOR2_NUM2257 (.ZN (N5950), .A1 (N5904), .A2 (N828));
      NOR2_X1 XNOR_NOR2_NUM2258 (.ZN (N5954), .A1 (N5858), .A2 (N5907));
      NOR2_X1 XNOR_NOR2_NUM2259 (.ZN (N5955), .A1 (N5907), .A2 (N876));
      NOR2_X1 XNOR_NOR2_NUM2260 (.ZN (N5956), .A1 (N5755), .A2 (N5907));
      NOR2_X1 XNOR_NOR2_NUM2261 (.ZN (N5959), .A1 (N5911), .A2 (N5912));
      NOR2_X1 XNOR_NOR2_NUM2262 (.ZN (N5962), .A1 (N5916), .A2 (N5913));
      NOR2_X1 XNOR_NOR2_NUM2263 (.ZN (N5966), .A1 (N5870), .A2 (N5919));
      NOR2_X1 XNOR_NOR2_NUM2264 (.ZN (N5967), .A1 (N5919), .A2 (N5867));
      NOR2_X1 XNOR_NOR2_NUM2265 (.ZN (N5968), .A1 (N5923), .A2 (N5924));
      NOR2_X1 XNOR_NOR2_NUM2266 (.ZN (N5971), .A1 (N5928), .A2 (N5929));
      NOR2_X1 XNOR_NOR2_NUM2267 (.ZN (N5972), .A1 (N5933), .A2 (N5934));
      NOR2_X1 XNOR_NOR2_NUM2268 (.ZN (N5975), .A1 (N5938), .A2 (N5935));
      NOR2_X1 XNOR_NOR2_NUM2269 (.ZN (N5979), .A1 (N5895), .A2 (N5941));
      NOR2_X1 XNOR_NOR2_NUM2270 (.ZN (N5980), .A1 (N5941), .A2 (N5892));
      NOR2_X1 XNOR_NOR2_NUM2271 (.ZN (N5981), .A1 (N5945), .A2 (N5946));
      NOR2_X1 XNOR_NOR2_NUM2272 (.ZN (N5984), .A1 (N5947), .A2 (N780));
      NOR2_X1 XNOR_NOR2_NUM2273 (.ZN (N5988), .A1 (N5904), .A2 (N5950));
      NOR2_X1 XNOR_NOR2_NUM2274 (.ZN (N5989), .A1 (N5950), .A2 (N828));
      NOR2_X1 XNOR_NOR2_NUM2275 (.ZN (N5990), .A1 (N5804), .A2 (N5950));
      NOR2_X1 XNOR_NOR2_NUM2276 (.ZN (N5993), .A1 (N5954), .A2 (N5955));
      NOR2_X1 XNOR_NOR2_NUM2277 (.ZN (N5996), .A1 (N5959), .A2 (N5956));
      NOR2_X1 XNOR_NOR2_NUM2278 (.ZN (N6000), .A1 (N5916), .A2 (N5962));
      NOR2_X1 XNOR_NOR2_NUM2279 (.ZN (N6001), .A1 (N5962), .A2 (N5913));
      NOR2_X1 XNOR_NOR2_NUM2280 (.ZN (N6002), .A1 (N5966), .A2 (N5967));
      NOR2_X1 XNOR_NOR2_NUM2281 (.ZN (N6005), .A1 (N5972), .A2 (N5930));
      NOR2_X1 XNOR_NOR2_NUM2282 (.ZN (N6009), .A1 (N5938), .A2 (N5975));
      NOR2_X1 XNOR_NOR2_NUM2283 (.ZN (N6010), .A1 (N5975), .A2 (N5935));
      NOR2_X1 XNOR_NOR2_NUM2284 (.ZN (N6011), .A1 (N5979), .A2 (N5980));
      NOR2_X1 XNOR_NOR2_NUM2285 (.ZN (N6014), .A1 (N5981), .A2 (N732));
      NOR2_X1 XNOR_NOR2_NUM2286 (.ZN (N6018), .A1 (N5947), .A2 (N5984));
      NOR2_X1 XNOR_NOR2_NUM2287 (.ZN (N6019), .A1 (N5984), .A2 (N780));
      NOR2_X1 XNOR_NOR2_NUM2288 (.ZN (N6020), .A1 (N5852), .A2 (N5984));
      NOR2_X1 XNOR_NOR2_NUM2289 (.ZN (N6023), .A1 (N5988), .A2 (N5989));
      NOR2_X1 XNOR_NOR2_NUM2290 (.ZN (N6026), .A1 (N5993), .A2 (N5990));
      NOR2_X1 XNOR_NOR2_NUM2291 (.ZN (N6030), .A1 (N5959), .A2 (N5996));
      NOR2_X1 XNOR_NOR2_NUM2292 (.ZN (N6031), .A1 (N5996), .A2 (N5956));
      NOR2_X1 XNOR_NOR2_NUM2293 (.ZN (N6032), .A1 (N6000), .A2 (N6001));
      NOR2_X1 XNOR_NOR2_NUM2294 (.ZN (N6035), .A1 (N5972), .A2 (N6005));
      NOR2_X1 XNOR_NOR2_NUM2295 (.ZN (N6036), .A1 (N6005), .A2 (N5930));
      NOR2_X1 XNOR_NOR2_NUM2296 (.ZN (N6037), .A1 (N6009), .A2 (N6010));
      NOR2_X1 XNOR_NOR2_NUM2297 (.ZN (N6040), .A1 (N6011), .A2 (N684));
      NOR2_X1 XNOR_NOR2_NUM2298 (.ZN (N6044), .A1 (N5981), .A2 (N6014));
      NOR2_X1 XNOR_NOR2_NUM2299 (.ZN (N6045), .A1 (N6014), .A2 (N732));
      NOR2_X1 XNOR_NOR2_NUM2300 (.ZN (N6046), .A1 (N5898), .A2 (N6014));
      NOR2_X1 XNOR_NOR2_NUM2301 (.ZN (N6049), .A1 (N6018), .A2 (N6019));
      NOR2_X1 XNOR_NOR2_NUM2302 (.ZN (N6052), .A1 (N6023), .A2 (N6020));
      NOR2_X1 XNOR_NOR2_NUM2303 (.ZN (N6056), .A1 (N5993), .A2 (N6026));
      NOR2_X1 XNOR_NOR2_NUM2304 (.ZN (N6057), .A1 (N6026), .A2 (N5990));
      NOR2_X1 XNOR_NOR2_NUM2305 (.ZN (N6058), .A1 (N6030), .A2 (N6031));
      NOR2_X1 XNOR_NOR2_NUM2306 (.ZN (N6061), .A1 (N6035), .A2 (N6036));
      NOR2_X1 XNOR_NOR2_NUM2307 (.ZN (N6064), .A1 (N6037), .A2 (N636));
      NOR2_X1 XNOR_NOR2_NUM2308 (.ZN (N6068), .A1 (N6011), .A2 (N6040));
      NOR2_X1 XNOR_NOR2_NUM2309 (.ZN (N6069), .A1 (N6040), .A2 (N684));
      NOR2_X1 XNOR_NOR2_NUM2310 (.ZN (N6070), .A1 (N5941), .A2 (N6040));
      NOR2_X1 XNOR_NOR2_NUM2311 (.ZN (N6073), .A1 (N6044), .A2 (N6045));
      NOR2_X1 XNOR_NOR2_NUM2312 (.ZN (N6076), .A1 (N6049), .A2 (N6046));
      NOR2_X1 XNOR_NOR2_NUM2313 (.ZN (N6080), .A1 (N6023), .A2 (N6052));
      NOR2_X1 XNOR_NOR2_NUM2314 (.ZN (N6081), .A1 (N6052), .A2 (N6020));
      NOR2_X1 XNOR_NOR2_NUM2315 (.ZN (N6082), .A1 (N6056), .A2 (N6057));
      NOR2_X1 XNOR_NOR2_NUM2316 (.ZN (N6085), .A1 (N6061), .A2 (N588));
      NOR2_X1 XNOR_NOR2_NUM2317 (.ZN (N6089), .A1 (N6037), .A2 (N6064));
      NOR2_X1 XNOR_NOR2_NUM2318 (.ZN (N6090), .A1 (N6064), .A2 (N636));
      NOR2_X1 XNOR_NOR2_NUM2319 (.ZN (N6091), .A1 (N5975), .A2 (N6064));
      NOR2_X1 XNOR_NOR2_NUM2320 (.ZN (N6094), .A1 (N6068), .A2 (N6069));
      NOR2_X1 XNOR_NOR2_NUM2321 (.ZN (N6097), .A1 (N6073), .A2 (N6070));
      NOR2_X1 XNOR_NOR2_NUM2322 (.ZN (N6101), .A1 (N6049), .A2 (N6076));
      NOR2_X1 XNOR_NOR2_NUM2323 (.ZN (N6102), .A1 (N6076), .A2 (N6046));
      NOR2_X1 XNOR_NOR2_NUM2324 (.ZN (N6103), .A1 (N6080), .A2 (N6081));
      NOR2_X1 XNOR_NOR2_NUM2325 (.ZN (N6106), .A1 (N6061), .A2 (N6085));
      NOR2_X1 XNOR_NOR2_NUM2326 (.ZN (N6107), .A1 (N6085), .A2 (N588));
      NOR2_X1 XNOR_NOR2_NUM2327 (.ZN (N6108), .A1 (N6005), .A2 (N6085));
      NOR2_X1 XNOR_NOR2_NUM2328 (.ZN (N6111), .A1 (N6089), .A2 (N6090));
      NOR2_X1 XNOR_NOR2_NUM2329 (.ZN (N6114), .A1 (N6094), .A2 (N6091));
      NOR2_X1 XNOR_NOR2_NUM2330 (.ZN (N6118), .A1 (N6073), .A2 (N6097));
      NOR2_X1 XNOR_NOR2_NUM2331 (.ZN (N6119), .A1 (N6097), .A2 (N6070));
      NOR2_X1 XNOR_NOR2_NUM2332 (.ZN (N6120), .A1 (N6101), .A2 (N6102));
      NOR2_X1 XNOR_NOR2_NUM2333 (.ZN (N6123), .A1 (N6106), .A2 (N6107));
      NOR2_X1 XNOR_NOR2_NUM2334 (.ZN (N6124), .A1 (N6111), .A2 (N6108));
      NOR2_X1 XNOR_NOR2_NUM2335 (.ZN (N6128), .A1 (N6094), .A2 (N6114));
      NOR2_X1 XNOR_NOR2_NUM2336 (.ZN (N6129), .A1 (N6114), .A2 (N6091));
      NOR2_X1 XNOR_NOR2_NUM2337 (.ZN (N6130), .A1 (N6118), .A2 (N6119));
      NOR2_X1 XNOR_NOR2_NUM2338 (.ZN (N6133), .A1 (N6111), .A2 (N6124));
      NOR2_X1 XNOR_NOR2_NUM2339 (.ZN (N6134), .A1 (N6124), .A2 (N6108));
      NOR2_X1 XNOR_NOR2_NUM2340 (.ZN (N6135), .A1 (N6128), .A2 (N6129));
      NOR2_X1 XNOR_NOR2_NUM2341 (.ZN (N6138), .A1 (N6133), .A2 (N6134));
      NOR2_X1 XNOR_NOT1_NUM2342 (.ZN (N6141), .A1 (N6138), .A2 (GND));
      NOR2_X1 XNOR_NOR2_NUM2343 (.ZN (N6145), .A1 (N6138), .A2 (N6141));
      NOR2_X1 XNOR_NOT1_NUM2344 (.ZN (N6146), .A1 (N6141), .A2 (GND));
      NOR2_X1 XNOR_NOR2_NUM2345 (.ZN (N6147), .A1 (N6124), .A2 (N6141));
      NOR2_X1 XNOR_NOR2_NUM2346 (.ZN (N6150), .A1 (N6145), .A2 (N6146));
      NOR2_X1 XNOR_NOR2_NUM2347 (.ZN (N6151), .A1 (N6135), .A2 (N6147));
      NOR2_X1 XNOR_NOR2_NUM2348 (.ZN (N6155), .A1 (N6135), .A2 (N6151));
      NOR2_X1 XNOR_NOR2_NUM2349 (.ZN (N6156), .A1 (N6151), .A2 (N6147));
      NOR2_X1 XNOR_NOR2_NUM2350 (.ZN (N6157), .A1 (N6114), .A2 (N6151));
      NOR2_X1 XNOR_NOR2_NUM2351 (.ZN (N6160), .A1 (N6155), .A2 (N6156));
      NOR2_X1 XNOR_NOR2_NUM2352 (.ZN (N6161), .A1 (N6130), .A2 (N6157));
      NOR2_X1 XNOR_NOR2_NUM2353 (.ZN (N6165), .A1 (N6130), .A2 (N6161));
      NOR2_X1 XNOR_NOR2_NUM2354 (.ZN (N6166), .A1 (N6161), .A2 (N6157));
      NOR2_X1 XNOR_NOR2_NUM2355 (.ZN (N6167), .A1 (N6097), .A2 (N6161));
      NOR2_X1 XNOR_NOR2_NUM2356 (.ZN (N6170), .A1 (N6165), .A2 (N6166));
      NOR2_X1 XNOR_NOR2_NUM2357 (.ZN (N6171), .A1 (N6120), .A2 (N6167));
      NOR2_X1 XNOR_NOR2_NUM2358 (.ZN (N6175), .A1 (N6120), .A2 (N6171));
      NOR2_X1 XNOR_NOR2_NUM2359 (.ZN (N6176), .A1 (N6171), .A2 (N6167));
      NOR2_X1 XNOR_NOR2_NUM2360 (.ZN (N6177), .A1 (N6076), .A2 (N6171));
      NOR2_X1 XNOR_NOR2_NUM2361 (.ZN (N6180), .A1 (N6175), .A2 (N6176));
      NOR2_X1 XNOR_NOR2_NUM2362 (.ZN (N6181), .A1 (N6103), .A2 (N6177));
      NOR2_X1 XNOR_NOR2_NUM2363 (.ZN (N6185), .A1 (N6103), .A2 (N6181));
      NOR2_X1 XNOR_NOR2_NUM2364 (.ZN (N6186), .A1 (N6181), .A2 (N6177));
      NOR2_X1 XNOR_NOR2_NUM2365 (.ZN (N6187), .A1 (N6052), .A2 (N6181));
      NOR2_X1 XNOR_NOR2_NUM2366 (.ZN (N6190), .A1 (N6185), .A2 (N6186));
      NOR2_X1 XNOR_NOR2_NUM2367 (.ZN (N6191), .A1 (N6082), .A2 (N6187));
      NOR2_X1 XNOR_NOR2_NUM2368 (.ZN (N6195), .A1 (N6082), .A2 (N6191));
      NOR2_X1 XNOR_NOR2_NUM2369 (.ZN (N6196), .A1 (N6191), .A2 (N6187));
      NOR2_X1 XNOR_NOR2_NUM2370 (.ZN (N6197), .A1 (N6026), .A2 (N6191));
      NOR2_X1 XNOR_NOR2_NUM2371 (.ZN (N6200), .A1 (N6195), .A2 (N6196));
      NOR2_X1 XNOR_NOR2_NUM2372 (.ZN (N6201), .A1 (N6058), .A2 (N6197));
      NOR2_X1 XNOR_NOR2_NUM2373 (.ZN (N6205), .A1 (N6058), .A2 (N6201));
      NOR2_X1 XNOR_NOR2_NUM2374 (.ZN (N6206), .A1 (N6201), .A2 (N6197));
      NOR2_X1 XNOR_NOR2_NUM2375 (.ZN (N6207), .A1 (N5996), .A2 (N6201));
      NOR2_X1 XNOR_NOR2_NUM2376 (.ZN (N6210), .A1 (N6205), .A2 (N6206));
      NOR2_X1 XNOR_NOR2_NUM2377 (.ZN (N6211), .A1 (N6032), .A2 (N6207));
      NOR2_X1 XNOR_NOR2_NUM2378 (.ZN (N6215), .A1 (N6032), .A2 (N6211));
      NOR2_X1 XNOR_NOR2_NUM2379 (.ZN (N6216), .A1 (N6211), .A2 (N6207));
      NOR2_X1 XNOR_NOR2_NUM2380 (.ZN (N6217), .A1 (N5962), .A2 (N6211));
      NOR2_X1 XNOR_NOR2_NUM2381 (.ZN (N6220), .A1 (N6215), .A2 (N6216));
      NOR2_X1 XNOR_NOR2_NUM2382 (.ZN (N6221), .A1 (N6002), .A2 (N6217));
      NOR2_X1 XNOR_NOR2_NUM2383 (.ZN (N6225), .A1 (N6002), .A2 (N6221));
      NOR2_X1 XNOR_NOR2_NUM2384 (.ZN (N6226), .A1 (N6221), .A2 (N6217));
      NOR2_X1 XNOR_NOR2_NUM2385 (.ZN (N6227), .A1 (N5919), .A2 (N6221));
      NOR2_X1 XNOR_NOR2_NUM2386 (.ZN (N6230), .A1 (N6225), .A2 (N6226));
      NOR2_X1 XNOR_NOR2_NUM2387 (.ZN (N6231), .A1 (N5968), .A2 (N6227));
      NOR2_X1 XNOR_NOR2_NUM2388 (.ZN (N6235), .A1 (N5968), .A2 (N6231));
      NOR2_X1 XNOR_NOR2_NUM2389 (.ZN (N6236), .A1 (N6231), .A2 (N6227));
      NOR2_X1 XNOR_NOR2_NUM2390 (.ZN (N6237), .A1 (N5873), .A2 (N6231));
      NOR2_X1 XNOR_NOR2_NUM2391 (.ZN (N6240), .A1 (N6235), .A2 (N6236));
      NOR2_X1 XNOR_NOR2_NUM2392 (.ZN (N6241), .A1 (N5925), .A2 (N6237));
      NOR2_X1 XNOR_NOR2_NUM2393 (.ZN (N6245), .A1 (N5925), .A2 (N6241));
      NOR2_X1 XNOR_NOR2_NUM2394 (.ZN (N6246), .A1 (N6241), .A2 (N6237));
      NOR2_X1 XNOR_NOR2_NUM2395 (.ZN (N6247), .A1 (N5825), .A2 (N6241));
      NOR2_X1 XNOR_NOR2_NUM2396 (.ZN (N6250), .A1 (N6245), .A2 (N6246));
      NOR2_X1 XNOR_NOR2_NUM2397 (.ZN (N6251), .A1 (N5879), .A2 (N6247));
      NOR2_X1 XNOR_NOR2_NUM2398 (.ZN (N6255), .A1 (N5879), .A2 (N6251));
      NOR2_X1 XNOR_NOR2_NUM2399 (.ZN (N6256), .A1 (N6251), .A2 (N6247));
      NOR2_X1 XNOR_NOR2_NUM2400 (.ZN (N6257), .A1 (N5776), .A2 (N6251));
      NOR2_X1 XNOR_NOR2_NUM2401 (.ZN (N6260), .A1 (N6255), .A2 (N6256));
      NOR2_X1 XNOR_NOR2_NUM2402 (.ZN (N6261), .A1 (N5831), .A2 (N6257));
      NOR2_X1 XNOR_NOR2_NUM2403 (.ZN (N6265), .A1 (N5831), .A2 (N6261));
      NOR2_X1 XNOR_NOR2_NUM2404 (.ZN (N6266), .A1 (N6261), .A2 (N6257));
      NOR2_X1 XNOR_NOR2_NUM2405 (.ZN (N6267), .A1 (N5721), .A2 (N6261));
      NOR2_X1 XNOR_NOR2_NUM2406 (.ZN (N6270), .A1 (N6265), .A2 (N6266));
      NOR2_X1 XNOR_NOR2_NUM2407 (.ZN (N6271), .A1 (N5782), .A2 (N6267));
      NOR2_X1 XNOR_NOR2_NUM2408 (.ZN (N6275), .A1 (N5782), .A2 (N6271));
      NOR2_X1 XNOR_NOR2_NUM2409 (.ZN (N6276), .A1 (N6271), .A2 (N6267));
      NOR2_X1 XNOR_NOR2_NUM2410 (.ZN (N6277), .A1 (N5666), .A2 (N6271));
      NOR2_X1 XNOR_NOR2_NUM2411 (.ZN (N6280), .A1 (N6275), .A2 (N6276));
      NOR2_X1 XNOR_NOR2_NUM2412 (.ZN (N6281), .A1 (N5727), .A2 (N6277));
      NOR2_X1 XNOR_NOR2_NUM2413 (.ZN (N6285), .A1 (N5727), .A2 (N6281));
      NOR2_X1 XNOR_NOR2_NUM2414 (.ZN (N6286), .A1 (N6281), .A2 (N6277));
      NOR2_X1 XNOR_NOR2_NUM2415 (.ZN (N6287), .A1 (N5602), .A2 (N6281));
      NOR2_X1 XNOR_NOR2_NUM2416 (.ZN (N6288), .A1 (N6285), .A2 (N6286));


      wire XNOR_1_1_N545_TERMINATION_OUT, XNOR_1_2_N545_TERMINATION_OUT;
      NOR2_X1 XNOR_1_1_N545_TERMINATION (.ZN (XNOR_1_1_N545_TERMINATION_OUT), .A1 (N545), .A2 (GND));
      NOR2_X1 XNOR_1_2_N545_TERMINATION (.ZN (N545_TERMINATION), .A1 (XNOR_1_1_N545_TERMINATION_OUT), .A2 (XNOR_1_2_N545_TERMINATION_OUT));

      wire XNOR_1_1_N1581_TERMINATION_OUT, XNOR_1_2_N1581_TERMINATION_OUT;
      NOR2_X1 XNOR_1_1_N1581_TERMINATION (.ZN (XNOR_1_1_N1581_TERMINATION_OUT), .A1 (N1581), .A2 (GND));
      NOR2_X1 XNOR_1_2_N1581_TERMINATION (.ZN (N1581_TERMINATION), .A1 (XNOR_1_1_N1581_TERMINATION_OUT), .A2 (XNOR_1_2_N1581_TERMINATION_OUT));

      wire XNOR_1_1_N1901_TERMINATION_OUT, XNOR_1_2_N1901_TERMINATION_OUT;
      NOR2_X1 XNOR_1_1_N1901_TERMINATION (.ZN (XNOR_1_1_N1901_TERMINATION_OUT), .A1 (N1901), .A2 (GND));
      NOR2_X1 XNOR_1_2_N1901_TERMINATION (.ZN (N1901_TERMINATION), .A1 (XNOR_1_1_N1901_TERMINATION_OUT), .A2 (XNOR_1_2_N1901_TERMINATION_OUT));

      wire XNOR_1_1_N2223_TERMINATION_OUT, XNOR_1_2_N2223_TERMINATION_OUT;
      NOR2_X1 XNOR_1_1_N2223_TERMINATION (.ZN (XNOR_1_1_N2223_TERMINATION_OUT), .A1 (N2223), .A2 (GND));
      NOR2_X1 XNOR_1_2_N2223_TERMINATION (.ZN (N2223_TERMINATION), .A1 (XNOR_1_1_N2223_TERMINATION_OUT), .A2 (XNOR_1_2_N2223_TERMINATION_OUT));

      wire XNOR_1_1_N2548_TERMINATION_OUT, XNOR_1_2_N2548_TERMINATION_OUT;
      NOR2_X1 XNOR_1_1_N2548_TERMINATION (.ZN (XNOR_1_1_N2548_TERMINATION_OUT), .A1 (N2548), .A2 (GND));
      NOR2_X1 XNOR_1_2_N2548_TERMINATION (.ZN (N2548_TERMINATION), .A1 (XNOR_1_1_N2548_TERMINATION_OUT), .A2 (XNOR_1_2_N2548_TERMINATION_OUT));

      wire XNOR_1_1_N2877_TERMINATION_OUT, XNOR_1_2_N2877_TERMINATION_OUT;
      NOR2_X1 XNOR_1_1_N2877_TERMINATION (.ZN (XNOR_1_1_N2877_TERMINATION_OUT), .A1 (N2877), .A2 (GND));
      NOR2_X1 XNOR_1_2_N2877_TERMINATION (.ZN (N2877_TERMINATION), .A1 (XNOR_1_1_N2877_TERMINATION_OUT), .A2 (XNOR_1_2_N2877_TERMINATION_OUT));

      wire XNOR_1_1_N3211_TERMINATION_OUT, XNOR_1_2_N3211_TERMINATION_OUT;
      NOR2_X1 XNOR_1_1_N3211_TERMINATION (.ZN (XNOR_1_1_N3211_TERMINATION_OUT), .A1 (N3211), .A2 (GND));
      NOR2_X1 XNOR_1_2_N3211_TERMINATION (.ZN (N3211_TERMINATION), .A1 (XNOR_1_1_N3211_TERMINATION_OUT), .A2 (XNOR_1_2_N3211_TERMINATION_OUT));

      wire XNOR_1_1_N3552_TERMINATION_OUT, XNOR_1_2_N3552_TERMINATION_OUT;
      NOR2_X1 XNOR_1_1_N3552_TERMINATION (.ZN (XNOR_1_1_N3552_TERMINATION_OUT), .A1 (N3552), .A2 (GND));
      NOR2_X1 XNOR_1_2_N3552_TERMINATION (.ZN (N3552_TERMINATION), .A1 (XNOR_1_1_N3552_TERMINATION_OUT), .A2 (XNOR_1_2_N3552_TERMINATION_OUT));

      wire XNOR_1_1_N3895_TERMINATION_OUT, XNOR_1_2_N3895_TERMINATION_OUT;
      NOR2_X1 XNOR_1_1_N3895_TERMINATION (.ZN (XNOR_1_1_N3895_TERMINATION_OUT), .A1 (N3895), .A2 (GND));
      NOR2_X1 XNOR_1_2_N3895_TERMINATION (.ZN (N3895_TERMINATION), .A1 (XNOR_1_1_N3895_TERMINATION_OUT), .A2 (XNOR_1_2_N3895_TERMINATION_OUT));

      wire XNOR_1_1_N4241_TERMINATION_OUT, XNOR_1_2_N4241_TERMINATION_OUT;
      NOR2_X1 XNOR_1_1_N4241_TERMINATION (.ZN (XNOR_1_1_N4241_TERMINATION_OUT), .A1 (N4241), .A2 (GND));
      NOR2_X1 XNOR_1_2_N4241_TERMINATION (.ZN (N4241_TERMINATION), .A1 (XNOR_1_1_N4241_TERMINATION_OUT), .A2 (XNOR_1_2_N4241_TERMINATION_OUT));

      wire XNOR_1_1_N4591_TERMINATION_OUT, XNOR_1_2_N4591_TERMINATION_OUT;
      NOR2_X1 XNOR_1_1_N4591_TERMINATION (.ZN (XNOR_1_1_N4591_TERMINATION_OUT), .A1 (N4591), .A2 (GND));
      NOR2_X1 XNOR_1_2_N4591_TERMINATION (.ZN (N4591_TERMINATION), .A1 (XNOR_1_1_N4591_TERMINATION_OUT), .A2 (XNOR_1_2_N4591_TERMINATION_OUT));

      wire XNOR_1_1_N4946_TERMINATION_OUT, XNOR_1_2_N4946_TERMINATION_OUT;
      NOR2_X1 XNOR_1_1_N4946_TERMINATION (.ZN (XNOR_1_1_N4946_TERMINATION_OUT), .A1 (N4946), .A2 (GND));
      NOR2_X1 XNOR_1_2_N4946_TERMINATION (.ZN (N4946_TERMINATION), .A1 (XNOR_1_1_N4946_TERMINATION_OUT), .A2 (XNOR_1_2_N4946_TERMINATION_OUT));

      wire XNOR_1_1_N5308_TERMINATION_OUT, XNOR_1_2_N5308_TERMINATION_OUT;
      NOR2_X1 XNOR_1_1_N5308_TERMINATION (.ZN (XNOR_1_1_N5308_TERMINATION_OUT), .A1 (N5308), .A2 (GND));
      NOR2_X1 XNOR_1_2_N5308_TERMINATION (.ZN (N5308_TERMINATION), .A1 (XNOR_1_1_N5308_TERMINATION_OUT), .A2 (XNOR_1_2_N5308_TERMINATION_OUT));

      wire XNOR_1_1_N5672_TERMINATION_OUT, XNOR_1_2_N5672_TERMINATION_OUT;
      NOR2_X1 XNOR_1_1_N5672_TERMINATION (.ZN (XNOR_1_1_N5672_TERMINATION_OUT), .A1 (N5672), .A2 (GND));
      NOR2_X1 XNOR_1_2_N5672_TERMINATION (.ZN (N5672_TERMINATION), .A1 (XNOR_1_1_N5672_TERMINATION_OUT), .A2 (XNOR_1_2_N5672_TERMINATION_OUT));

      wire XNOR_1_1_N5971_TERMINATION_OUT, XNOR_1_2_N5971_TERMINATION_OUT;
      NOR2_X1 XNOR_1_1_N5971_TERMINATION (.ZN (XNOR_1_1_N5971_TERMINATION_OUT), .A1 (N5971), .A2 (GND));
      NOR2_X1 XNOR_1_2_N5971_TERMINATION (.ZN (N5971_TERMINATION), .A1 (XNOR_1_1_N5971_TERMINATION_OUT), .A2 (XNOR_1_2_N5971_TERMINATION_OUT));

      wire XNOR_1_1_N6123_TERMINATION_OUT, XNOR_1_2_N6123_TERMINATION_OUT;
      NOR2_X1 XNOR_1_1_N6123_TERMINATION (.ZN (XNOR_1_1_N6123_TERMINATION_OUT), .A1 (N6123), .A2 (GND));
      NOR2_X1 XNOR_1_2_N6123_TERMINATION (.ZN (N6123_TERMINATION), .A1 (XNOR_1_1_N6123_TERMINATION_OUT), .A2 (XNOR_1_2_N6123_TERMINATION_OUT));

      wire XNOR_1_1_N6150_TERMINATION_OUT, XNOR_1_2_N6150_TERMINATION_OUT;
      NOR2_X1 XNOR_1_1_N6150_TERMINATION (.ZN (XNOR_1_1_N6150_TERMINATION_OUT), .A1 (N6150), .A2 (GND));
      NOR2_X1 XNOR_1_2_N6150_TERMINATION (.ZN (N6150_TERMINATION), .A1 (XNOR_1_1_N6150_TERMINATION_OUT), .A2 (XNOR_1_2_N6150_TERMINATION_OUT));

      wire XNOR_1_1_N6160_TERMINATION_OUT, XNOR_1_2_N6160_TERMINATION_OUT;
      NOR2_X1 XNOR_1_1_N6160_TERMINATION (.ZN (XNOR_1_1_N6160_TERMINATION_OUT), .A1 (N6160), .A2 (GND));
      NOR2_X1 XNOR_1_2_N6160_TERMINATION (.ZN (N6160_TERMINATION), .A1 (XNOR_1_1_N6160_TERMINATION_OUT), .A2 (XNOR_1_2_N6160_TERMINATION_OUT));

      wire XNOR_1_1_N6170_TERMINATION_OUT, XNOR_1_2_N6170_TERMINATION_OUT;
      NOR2_X1 XNOR_1_1_N6170_TERMINATION (.ZN (XNOR_1_1_N6170_TERMINATION_OUT), .A1 (N6170), .A2 (GND));
      NOR2_X1 XNOR_1_2_N6170_TERMINATION (.ZN (N6170_TERMINATION), .A1 (XNOR_1_1_N6170_TERMINATION_OUT), .A2 (XNOR_1_2_N6170_TERMINATION_OUT));

      wire XNOR_1_1_N6180_TERMINATION_OUT, XNOR_1_2_N6180_TERMINATION_OUT;
      NOR2_X1 XNOR_1_1_N6180_TERMINATION (.ZN (XNOR_1_1_N6180_TERMINATION_OUT), .A1 (N6180), .A2 (GND));
      NOR2_X1 XNOR_1_2_N6180_TERMINATION (.ZN (N6180_TERMINATION), .A1 (XNOR_1_1_N6180_TERMINATION_OUT), .A2 (XNOR_1_2_N6180_TERMINATION_OUT));

      wire XNOR_1_1_N6190_TERMINATION_OUT, XNOR_1_2_N6190_TERMINATION_OUT;
      NOR2_X1 XNOR_1_1_N6190_TERMINATION (.ZN (XNOR_1_1_N6190_TERMINATION_OUT), .A1 (N6190), .A2 (GND));
      NOR2_X1 XNOR_1_2_N6190_TERMINATION (.ZN (N6190_TERMINATION), .A1 (XNOR_1_1_N6190_TERMINATION_OUT), .A2 (XNOR_1_2_N6190_TERMINATION_OUT));

      wire XNOR_1_1_N6200_TERMINATION_OUT, XNOR_1_2_N6200_TERMINATION_OUT;
      NOR2_X1 XNOR_1_1_N6200_TERMINATION (.ZN (XNOR_1_1_N6200_TERMINATION_OUT), .A1 (N6200), .A2 (GND));
      NOR2_X1 XNOR_1_2_N6200_TERMINATION (.ZN (N6200_TERMINATION), .A1 (XNOR_1_1_N6200_TERMINATION_OUT), .A2 (XNOR_1_2_N6200_TERMINATION_OUT));

      wire XNOR_1_1_N6210_TERMINATION_OUT, XNOR_1_2_N6210_TERMINATION_OUT;
      NOR2_X1 XNOR_1_1_N6210_TERMINATION (.ZN (XNOR_1_1_N6210_TERMINATION_OUT), .A1 (N6210), .A2 (GND));
      NOR2_X1 XNOR_1_2_N6210_TERMINATION (.ZN (N6210_TERMINATION), .A1 (XNOR_1_1_N6210_TERMINATION_OUT), .A2 (XNOR_1_2_N6210_TERMINATION_OUT));

      wire XNOR_1_1_N6220_TERMINATION_OUT, XNOR_1_2_N6220_TERMINATION_OUT;
      NOR2_X1 XNOR_1_1_N6220_TERMINATION (.ZN (XNOR_1_1_N6220_TERMINATION_OUT), .A1 (N6220), .A2 (GND));
      NOR2_X1 XNOR_1_2_N6220_TERMINATION (.ZN (N6220_TERMINATION), .A1 (XNOR_1_1_N6220_TERMINATION_OUT), .A2 (XNOR_1_2_N6220_TERMINATION_OUT));

      wire XNOR_1_1_N6230_TERMINATION_OUT, XNOR_1_2_N6230_TERMINATION_OUT;
      NOR2_X1 XNOR_1_1_N6230_TERMINATION (.ZN (XNOR_1_1_N6230_TERMINATION_OUT), .A1 (N6230), .A2 (GND));
      NOR2_X1 XNOR_1_2_N6230_TERMINATION (.ZN (N6230_TERMINATION), .A1 (XNOR_1_1_N6230_TERMINATION_OUT), .A2 (XNOR_1_2_N6230_TERMINATION_OUT));

      wire XNOR_1_1_N6240_TERMINATION_OUT, XNOR_1_2_N6240_TERMINATION_OUT;
      NOR2_X1 XNOR_1_1_N6240_TERMINATION (.ZN (XNOR_1_1_N6240_TERMINATION_OUT), .A1 (N6240), .A2 (GND));
      NOR2_X1 XNOR_1_2_N6240_TERMINATION (.ZN (N6240_TERMINATION), .A1 (XNOR_1_1_N6240_TERMINATION_OUT), .A2 (XNOR_1_2_N6240_TERMINATION_OUT));

      wire XNOR_1_1_N6250_TERMINATION_OUT, XNOR_1_2_N6250_TERMINATION_OUT;
      NOR2_X1 XNOR_1_1_N6250_TERMINATION (.ZN (XNOR_1_1_N6250_TERMINATION_OUT), .A1 (N6250), .A2 (GND));
      NOR2_X1 XNOR_1_2_N6250_TERMINATION (.ZN (N6250_TERMINATION), .A1 (XNOR_1_1_N6250_TERMINATION_OUT), .A2 (XNOR_1_2_N6250_TERMINATION_OUT));

      wire XNOR_1_1_N6260_TERMINATION_OUT, XNOR_1_2_N6260_TERMINATION_OUT;
      NOR2_X1 XNOR_1_1_N6260_TERMINATION (.ZN (XNOR_1_1_N6260_TERMINATION_OUT), .A1 (N6260), .A2 (GND));
      NOR2_X1 XNOR_1_2_N6260_TERMINATION (.ZN (N6260_TERMINATION), .A1 (XNOR_1_1_N6260_TERMINATION_OUT), .A2 (XNOR_1_2_N6260_TERMINATION_OUT));

      wire XNOR_1_1_N6270_TERMINATION_OUT, XNOR_1_2_N6270_TERMINATION_OUT;
      NOR2_X1 XNOR_1_1_N6270_TERMINATION (.ZN (XNOR_1_1_N6270_TERMINATION_OUT), .A1 (N6270), .A2 (GND));
      NOR2_X1 XNOR_1_2_N6270_TERMINATION (.ZN (N6270_TERMINATION), .A1 (XNOR_1_1_N6270_TERMINATION_OUT), .A2 (XNOR_1_2_N6270_TERMINATION_OUT));

      wire XNOR_1_1_N6280_TERMINATION_OUT, XNOR_1_2_N6280_TERMINATION_OUT;
      NOR2_X1 XNOR_1_1_N6280_TERMINATION (.ZN (XNOR_1_1_N6280_TERMINATION_OUT), .A1 (N6280), .A2 (GND));
      NOR2_X1 XNOR_1_2_N6280_TERMINATION (.ZN (N6280_TERMINATION), .A1 (XNOR_1_1_N6280_TERMINATION_OUT), .A2 (XNOR_1_2_N6280_TERMINATION_OUT));

      wire XNOR_1_1_N6287_TERMINATION_OUT, XNOR_1_2_N6287_TERMINATION_OUT;
      NOR2_X1 XNOR_1_1_N6287_TERMINATION (.ZN (XNOR_1_1_N6287_TERMINATION_OUT), .A1 (N6287), .A2 (GND));
      NOR2_X1 XNOR_1_2_N6287_TERMINATION (.ZN (N6287_TERMINATION), .A1 (XNOR_1_1_N6287_TERMINATION_OUT), .A2 (XNOR_1_2_N6287_TERMINATION_OUT));

      wire XNOR_1_1_N6288_TERMINATION_OUT, XNOR_1_2_N6288_TERMINATION_OUT;
      NOR2_X1 XNOR_1_1_N6288_TERMINATION (.ZN (XNOR_1_1_N6288_TERMINATION_OUT), .A1 (N6288), .A2 (GND));
      NOR2_X1 XNOR_1_2_N6288_TERMINATION (.ZN (N6288_TERMINATION), .A1 (XNOR_1_1_N6288_TERMINATION_OUT), .A2 (XNOR_1_2_N6288_TERMINATION_OUT));




endmodule
module c1355_NOR_template (N1_PWL,N8_PWL,N15_PWL,N22_PWL,N29_PWL,N36_PWL,N43_PWL,N50_PWL,N57_PWL,N64_PWL,N71_PWL,N78_PWL,N85_PWL,N92_PWL,N99_PWL,N106_PWL,N113_PWL,N120_PWL,N127_PWL,N134_PWL,
            N141_PWL,N148_PWL,N155_PWL,N162_PWL,N169_PWL,N176_PWL,N183_PWL,N190_PWL,N197_PWL,N204_PWL,N211_PWL,N218_PWL,N225_PWL,N226_PWL,N227_PWL,N228_PWL,N229_PWL,
            N230_PWL,N231_PWL,N232_PWL,N233_PWL,
            N1324_TERMINATION,N1325_TERMINATION,N1326_TERMINATION,N1327_TERMINATION,N1328_TERMINATION,N1329_TERMINATION,N1330_TERMINATION,N1331_TERMINATION,N1332_TERMINATION,N1333_TERMINATION,N1334_TERMINATION,N1335_TERMINATION,N1336_TERMINATION,N1337_TERMINATION,
            N1338_TERMINATION,N1339_TERMINATION,N1340_TERMINATION,N1341_TERMINATION,N1342_TERMINATION,N1343_TERMINATION,N1344_TERMINATION,N1345_TERMINATION,N1346_TERMINATION,N1347_TERMINATION,N1348_TERMINATION,N1349_TERMINATION,N1350_TERMINATION,N1351_TERMINATION,
            N1352_TERMINATION,N1353_TERMINATION,N1354_TERMINATION,N1355_TERMINATION);

      input N1_PWL,N8_PWL,N15_PWL,N22_PWL,N29_PWL,N36_PWL,N43_PWL,N50_PWL,N57_PWL,N64_PWL,N71_PWL,N78_PWL,N85_PWL,N92_PWL,N99_PWL,N106_PWL,N113_PWL,N120_PWL,N127_PWL,N134_PWL,
            N141_PWL,N148_PWL,N155_PWL,N162_PWL,N169_PWL,N176_PWL,N183_PWL,N190_PWL,N197_PWL,N204_PWL,N211_PWL,N218_PWL,N225_PWL,N226_PWL,N227_PWL,N228_PWL,N229_PWL,
            N230_PWL,N231_PWL,N232_PWL,N233_PWL;

      output N1324_TERMINATION,N1325_TERMINATION,N1326_TERMINATION,N1327_TERMINATION,N1328_TERMINATION,N1329_TERMINATION,N1330_TERMINATION,N1331_TERMINATION,N1332_TERMINATION,N1333_TERMINATION,N1334_TERMINATION,N1335_TERMINATION,N1336_TERMINATION,N1337_TERMINATION,
            N1338_TERMINATION,N1339_TERMINATION,N1340_TERMINATION,N1341_TERMINATION,N1342_TERMINATION,N1343_TERMINATION,N1344_TERMINATION,N1345_TERMINATION,N1346_TERMINATION,N1347_TERMINATION,N1348_TERMINATION,N1349_TERMINATION,N1350_TERMINATION,N1351_TERMINATION,
            N1352_TERMINATION,N1353_TERMINATION,N1354_TERMINATION,N1355_TERMINATION;


      wire GND = 1'b0;
      wire XNOR_1_1_N1_PULSESHAPING_OUT, XNOR_1_2_N1_PULSESHAPING_OUT, XNOR_1_3_N1_PULSESHAPING_OUT, XNOR_1_4_N1_PULSESHAPING_OUT, XNOR_1_5_N1_PULSESHAPING_OUT, XNOR_1_6_N1_PULSESHAPING_OUT;
      NOR2_X1 XNOR_1_1_N1_PULSESHAPING (.ZN (XNOR_1_1_N1_PULSESHAPING_OUT), .A1 (N1_PWL), .A2 (GND));
      NOR2_X1 XNOR_1_2_N1_PULSESHAPING (.ZN (XNOR_1_2_N1_PULSESHAPING_OUT), .A1 (XNOR_1_1_N1_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_3_N1_PULSESHAPING (.ZN (XNOR_1_3_N1_PULSESHAPING_OUT), .A1 (XNOR_1_2_N1_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_4_N1_PULSESHAPING (.ZN (XNOR_1_4_N1_PULSESHAPING_OUT), .A1 (XNOR_1_3_N1_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_5_N1_PULSESHAPING (.ZN (XNOR_1_5_N1_PULSESHAPING_OUT), .A1 (XNOR_1_4_N1_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_6_N1_PULSESHAPING (.ZN (XNOR_1_6_N1_PULSESHAPING_OUT), .A1 (XNOR_1_5_N1_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_7_N1_PULSESHAPING (.ZN (N1), .A1 (XNOR_1_6_N1_PULSESHAPING_OUT), .A2 (GND));

      wire XNOR_1_1_N8_PULSESHAPING_OUT, XNOR_1_2_N8_PULSESHAPING_OUT, XNOR_1_3_N8_PULSESHAPING_OUT, XNOR_1_4_N8_PULSESHAPING_OUT, XNOR_1_5_N8_PULSESHAPING_OUT, XNOR_1_6_N8_PULSESHAPING_OUT;
      NOR2_X1 XNOR_1_1_N8_PULSESHAPING (.ZN (XNOR_1_1_N8_PULSESHAPING_OUT), .A1 (N8_PWL), .A2 (GND));
      NOR2_X1 XNOR_1_2_N8_PULSESHAPING (.ZN (XNOR_1_2_N8_PULSESHAPING_OUT), .A1 (XNOR_1_1_N8_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_3_N8_PULSESHAPING (.ZN (XNOR_1_3_N8_PULSESHAPING_OUT), .A1 (XNOR_1_2_N8_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_4_N8_PULSESHAPING (.ZN (XNOR_1_4_N8_PULSESHAPING_OUT), .A1 (XNOR_1_3_N8_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_5_N8_PULSESHAPING (.ZN (XNOR_1_5_N8_PULSESHAPING_OUT), .A1 (XNOR_1_4_N8_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_6_N8_PULSESHAPING (.ZN (XNOR_1_6_N8_PULSESHAPING_OUT), .A1 (XNOR_1_5_N8_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_7_N8_PULSESHAPING (.ZN (N8), .A1 (XNOR_1_6_N8_PULSESHAPING_OUT), .A2 (GND));

      wire XNOR_1_1_N15_PULSESHAPING_OUT, XNOR_1_2_N15_PULSESHAPING_OUT, XNOR_1_3_N15_PULSESHAPING_OUT, XNOR_1_4_N15_PULSESHAPING_OUT, XNOR_1_5_N15_PULSESHAPING_OUT, XNOR_1_6_N15_PULSESHAPING_OUT;
      NOR2_X1 XNOR_1_1_N15_PULSESHAPING (.ZN (XNOR_1_1_N15_PULSESHAPING_OUT), .A1 (N15_PWL), .A2 (GND));
      NOR2_X1 XNOR_1_2_N15_PULSESHAPING (.ZN (XNOR_1_2_N15_PULSESHAPING_OUT), .A1 (XNOR_1_1_N15_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_3_N15_PULSESHAPING (.ZN (XNOR_1_3_N15_PULSESHAPING_OUT), .A1 (XNOR_1_2_N15_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_4_N15_PULSESHAPING (.ZN (XNOR_1_4_N15_PULSESHAPING_OUT), .A1 (XNOR_1_3_N15_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_5_N15_PULSESHAPING (.ZN (XNOR_1_5_N15_PULSESHAPING_OUT), .A1 (XNOR_1_4_N15_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_6_N15_PULSESHAPING (.ZN (XNOR_1_6_N15_PULSESHAPING_OUT), .A1 (XNOR_1_5_N15_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_7_N15_PULSESHAPING (.ZN (N15), .A1 (XNOR_1_6_N15_PULSESHAPING_OUT), .A2 (GND));

      wire XNOR_1_1_N22_PULSESHAPING_OUT, XNOR_1_2_N22_PULSESHAPING_OUT, XNOR_1_3_N22_PULSESHAPING_OUT, XNOR_1_4_N22_PULSESHAPING_OUT, XNOR_1_5_N22_PULSESHAPING_OUT, XNOR_1_6_N22_PULSESHAPING_OUT;
      NOR2_X1 XNOR_1_1_N22_PULSESHAPING (.ZN (XNOR_1_1_N22_PULSESHAPING_OUT), .A1 (N22_PWL), .A2 (GND));
      NOR2_X1 XNOR_1_2_N22_PULSESHAPING (.ZN (XNOR_1_2_N22_PULSESHAPING_OUT), .A1 (XNOR_1_1_N22_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_3_N22_PULSESHAPING (.ZN (XNOR_1_3_N22_PULSESHAPING_OUT), .A1 (XNOR_1_2_N22_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_4_N22_PULSESHAPING (.ZN (XNOR_1_4_N22_PULSESHAPING_OUT), .A1 (XNOR_1_3_N22_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_5_N22_PULSESHAPING (.ZN (XNOR_1_5_N22_PULSESHAPING_OUT), .A1 (XNOR_1_4_N22_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_6_N22_PULSESHAPING (.ZN (XNOR_1_6_N22_PULSESHAPING_OUT), .A1 (XNOR_1_5_N22_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_7_N22_PULSESHAPING (.ZN (N22), .A1 (XNOR_1_6_N22_PULSESHAPING_OUT), .A2 (GND));

      wire XNOR_1_1_N29_PULSESHAPING_OUT, XNOR_1_2_N29_PULSESHAPING_OUT, XNOR_1_3_N29_PULSESHAPING_OUT, XNOR_1_4_N29_PULSESHAPING_OUT, XNOR_1_5_N29_PULSESHAPING_OUT, XNOR_1_6_N29_PULSESHAPING_OUT;
      NOR2_X1 XNOR_1_1_N29_PULSESHAPING (.ZN (XNOR_1_1_N29_PULSESHAPING_OUT), .A1 (N29_PWL), .A2 (GND));
      NOR2_X1 XNOR_1_2_N29_PULSESHAPING (.ZN (XNOR_1_2_N29_PULSESHAPING_OUT), .A1 (XNOR_1_1_N29_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_3_N29_PULSESHAPING (.ZN (XNOR_1_3_N29_PULSESHAPING_OUT), .A1 (XNOR_1_2_N29_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_4_N29_PULSESHAPING (.ZN (XNOR_1_4_N29_PULSESHAPING_OUT), .A1 (XNOR_1_3_N29_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_5_N29_PULSESHAPING (.ZN (XNOR_1_5_N29_PULSESHAPING_OUT), .A1 (XNOR_1_4_N29_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_6_N29_PULSESHAPING (.ZN (XNOR_1_6_N29_PULSESHAPING_OUT), .A1 (XNOR_1_5_N29_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_7_N29_PULSESHAPING (.ZN (N29), .A1 (XNOR_1_6_N29_PULSESHAPING_OUT), .A2 (GND));

      wire XNOR_1_1_N36_PULSESHAPING_OUT, XNOR_1_2_N36_PULSESHAPING_OUT, XNOR_1_3_N36_PULSESHAPING_OUT, XNOR_1_4_N36_PULSESHAPING_OUT, XNOR_1_5_N36_PULSESHAPING_OUT, XNOR_1_6_N36_PULSESHAPING_OUT;
      NOR2_X1 XNOR_1_1_N36_PULSESHAPING (.ZN (XNOR_1_1_N36_PULSESHAPING_OUT), .A1 (N36_PWL), .A2 (GND));
      NOR2_X1 XNOR_1_2_N36_PULSESHAPING (.ZN (XNOR_1_2_N36_PULSESHAPING_OUT), .A1 (XNOR_1_1_N36_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_3_N36_PULSESHAPING (.ZN (XNOR_1_3_N36_PULSESHAPING_OUT), .A1 (XNOR_1_2_N36_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_4_N36_PULSESHAPING (.ZN (XNOR_1_4_N36_PULSESHAPING_OUT), .A1 (XNOR_1_3_N36_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_5_N36_PULSESHAPING (.ZN (XNOR_1_5_N36_PULSESHAPING_OUT), .A1 (XNOR_1_4_N36_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_6_N36_PULSESHAPING (.ZN (XNOR_1_6_N36_PULSESHAPING_OUT), .A1 (XNOR_1_5_N36_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_7_N36_PULSESHAPING (.ZN (N36), .A1 (XNOR_1_6_N36_PULSESHAPING_OUT), .A2 (GND));

      wire XNOR_1_1_N43_PULSESHAPING_OUT, XNOR_1_2_N43_PULSESHAPING_OUT, XNOR_1_3_N43_PULSESHAPING_OUT, XNOR_1_4_N43_PULSESHAPING_OUT, XNOR_1_5_N43_PULSESHAPING_OUT, XNOR_1_6_N43_PULSESHAPING_OUT;
      NOR2_X1 XNOR_1_1_N43_PULSESHAPING (.ZN (XNOR_1_1_N43_PULSESHAPING_OUT), .A1 (N43_PWL), .A2 (GND));
      NOR2_X1 XNOR_1_2_N43_PULSESHAPING (.ZN (XNOR_1_2_N43_PULSESHAPING_OUT), .A1 (XNOR_1_1_N43_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_3_N43_PULSESHAPING (.ZN (XNOR_1_3_N43_PULSESHAPING_OUT), .A1 (XNOR_1_2_N43_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_4_N43_PULSESHAPING (.ZN (XNOR_1_4_N43_PULSESHAPING_OUT), .A1 (XNOR_1_3_N43_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_5_N43_PULSESHAPING (.ZN (XNOR_1_5_N43_PULSESHAPING_OUT), .A1 (XNOR_1_4_N43_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_6_N43_PULSESHAPING (.ZN (XNOR_1_6_N43_PULSESHAPING_OUT), .A1 (XNOR_1_5_N43_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_7_N43_PULSESHAPING (.ZN (N43), .A1 (XNOR_1_6_N43_PULSESHAPING_OUT), .A2 (GND));

      wire XNOR_1_1_N50_PULSESHAPING_OUT, XNOR_1_2_N50_PULSESHAPING_OUT, XNOR_1_3_N50_PULSESHAPING_OUT, XNOR_1_4_N50_PULSESHAPING_OUT, XNOR_1_5_N50_PULSESHAPING_OUT, XNOR_1_6_N50_PULSESHAPING_OUT;
      NOR2_X1 XNOR_1_1_N50_PULSESHAPING (.ZN (XNOR_1_1_N50_PULSESHAPING_OUT), .A1 (N50_PWL), .A2 (GND));
      NOR2_X1 XNOR_1_2_N50_PULSESHAPING (.ZN (XNOR_1_2_N50_PULSESHAPING_OUT), .A1 (XNOR_1_1_N50_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_3_N50_PULSESHAPING (.ZN (XNOR_1_3_N50_PULSESHAPING_OUT), .A1 (XNOR_1_2_N50_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_4_N50_PULSESHAPING (.ZN (XNOR_1_4_N50_PULSESHAPING_OUT), .A1 (XNOR_1_3_N50_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_5_N50_PULSESHAPING (.ZN (XNOR_1_5_N50_PULSESHAPING_OUT), .A1 (XNOR_1_4_N50_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_6_N50_PULSESHAPING (.ZN (XNOR_1_6_N50_PULSESHAPING_OUT), .A1 (XNOR_1_5_N50_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_7_N50_PULSESHAPING (.ZN (N50), .A1 (XNOR_1_6_N50_PULSESHAPING_OUT), .A2 (GND));

      wire XNOR_1_1_N57_PULSESHAPING_OUT, XNOR_1_2_N57_PULSESHAPING_OUT, XNOR_1_3_N57_PULSESHAPING_OUT, XNOR_1_4_N57_PULSESHAPING_OUT, XNOR_1_5_N57_PULSESHAPING_OUT, XNOR_1_6_N57_PULSESHAPING_OUT;
      NOR2_X1 XNOR_1_1_N57_PULSESHAPING (.ZN (XNOR_1_1_N57_PULSESHAPING_OUT), .A1 (N57_PWL), .A2 (GND));
      NOR2_X1 XNOR_1_2_N57_PULSESHAPING (.ZN (XNOR_1_2_N57_PULSESHAPING_OUT), .A1 (XNOR_1_1_N57_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_3_N57_PULSESHAPING (.ZN (XNOR_1_3_N57_PULSESHAPING_OUT), .A1 (XNOR_1_2_N57_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_4_N57_PULSESHAPING (.ZN (XNOR_1_4_N57_PULSESHAPING_OUT), .A1 (XNOR_1_3_N57_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_5_N57_PULSESHAPING (.ZN (XNOR_1_5_N57_PULSESHAPING_OUT), .A1 (XNOR_1_4_N57_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_6_N57_PULSESHAPING (.ZN (XNOR_1_6_N57_PULSESHAPING_OUT), .A1 (XNOR_1_5_N57_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_7_N57_PULSESHAPING (.ZN (N57), .A1 (XNOR_1_6_N57_PULSESHAPING_OUT), .A2 (GND));

      wire XNOR_1_1_N64_PULSESHAPING_OUT, XNOR_1_2_N64_PULSESHAPING_OUT, XNOR_1_3_N64_PULSESHAPING_OUT, XNOR_1_4_N64_PULSESHAPING_OUT, XNOR_1_5_N64_PULSESHAPING_OUT, XNOR_1_6_N64_PULSESHAPING_OUT;
      NOR2_X1 XNOR_1_1_N64_PULSESHAPING (.ZN (XNOR_1_1_N64_PULSESHAPING_OUT), .A1 (N64_PWL), .A2 (GND));
      NOR2_X1 XNOR_1_2_N64_PULSESHAPING (.ZN (XNOR_1_2_N64_PULSESHAPING_OUT), .A1 (XNOR_1_1_N64_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_3_N64_PULSESHAPING (.ZN (XNOR_1_3_N64_PULSESHAPING_OUT), .A1 (XNOR_1_2_N64_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_4_N64_PULSESHAPING (.ZN (XNOR_1_4_N64_PULSESHAPING_OUT), .A1 (XNOR_1_3_N64_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_5_N64_PULSESHAPING (.ZN (XNOR_1_5_N64_PULSESHAPING_OUT), .A1 (XNOR_1_4_N64_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_6_N64_PULSESHAPING (.ZN (XNOR_1_6_N64_PULSESHAPING_OUT), .A1 (XNOR_1_5_N64_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_7_N64_PULSESHAPING (.ZN (N64), .A1 (XNOR_1_6_N64_PULSESHAPING_OUT), .A2 (GND));

      wire XNOR_1_1_N71_PULSESHAPING_OUT, XNOR_1_2_N71_PULSESHAPING_OUT, XNOR_1_3_N71_PULSESHAPING_OUT, XNOR_1_4_N71_PULSESHAPING_OUT, XNOR_1_5_N71_PULSESHAPING_OUT, XNOR_1_6_N71_PULSESHAPING_OUT;
      NOR2_X1 XNOR_1_1_N71_PULSESHAPING (.ZN (XNOR_1_1_N71_PULSESHAPING_OUT), .A1 (N71_PWL), .A2 (GND));
      NOR2_X1 XNOR_1_2_N71_PULSESHAPING (.ZN (XNOR_1_2_N71_PULSESHAPING_OUT), .A1 (XNOR_1_1_N71_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_3_N71_PULSESHAPING (.ZN (XNOR_1_3_N71_PULSESHAPING_OUT), .A1 (XNOR_1_2_N71_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_4_N71_PULSESHAPING (.ZN (XNOR_1_4_N71_PULSESHAPING_OUT), .A1 (XNOR_1_3_N71_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_5_N71_PULSESHAPING (.ZN (XNOR_1_5_N71_PULSESHAPING_OUT), .A1 (XNOR_1_4_N71_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_6_N71_PULSESHAPING (.ZN (XNOR_1_6_N71_PULSESHAPING_OUT), .A1 (XNOR_1_5_N71_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_7_N71_PULSESHAPING (.ZN (N71), .A1 (XNOR_1_6_N71_PULSESHAPING_OUT), .A2 (GND));

      wire XNOR_1_1_N78_PULSESHAPING_OUT, XNOR_1_2_N78_PULSESHAPING_OUT, XNOR_1_3_N78_PULSESHAPING_OUT, XNOR_1_4_N78_PULSESHAPING_OUT, XNOR_1_5_N78_PULSESHAPING_OUT, XNOR_1_6_N78_PULSESHAPING_OUT;
      NOR2_X1 XNOR_1_1_N78_PULSESHAPING (.ZN (XNOR_1_1_N78_PULSESHAPING_OUT), .A1 (N78_PWL), .A2 (GND));
      NOR2_X1 XNOR_1_2_N78_PULSESHAPING (.ZN (XNOR_1_2_N78_PULSESHAPING_OUT), .A1 (XNOR_1_1_N78_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_3_N78_PULSESHAPING (.ZN (XNOR_1_3_N78_PULSESHAPING_OUT), .A1 (XNOR_1_2_N78_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_4_N78_PULSESHAPING (.ZN (XNOR_1_4_N78_PULSESHAPING_OUT), .A1 (XNOR_1_3_N78_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_5_N78_PULSESHAPING (.ZN (XNOR_1_5_N78_PULSESHAPING_OUT), .A1 (XNOR_1_4_N78_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_6_N78_PULSESHAPING (.ZN (XNOR_1_6_N78_PULSESHAPING_OUT), .A1 (XNOR_1_5_N78_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_7_N78_PULSESHAPING (.ZN (N78), .A1 (XNOR_1_6_N78_PULSESHAPING_OUT), .A2 (GND));

      wire XNOR_1_1_N85_PULSESHAPING_OUT, XNOR_1_2_N85_PULSESHAPING_OUT, XNOR_1_3_N85_PULSESHAPING_OUT, XNOR_1_4_N85_PULSESHAPING_OUT, XNOR_1_5_N85_PULSESHAPING_OUT, XNOR_1_6_N85_PULSESHAPING_OUT;
      NOR2_X1 XNOR_1_1_N85_PULSESHAPING (.ZN (XNOR_1_1_N85_PULSESHAPING_OUT), .A1 (N85_PWL), .A2 (GND));
      NOR2_X1 XNOR_1_2_N85_PULSESHAPING (.ZN (XNOR_1_2_N85_PULSESHAPING_OUT), .A1 (XNOR_1_1_N85_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_3_N85_PULSESHAPING (.ZN (XNOR_1_3_N85_PULSESHAPING_OUT), .A1 (XNOR_1_2_N85_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_4_N85_PULSESHAPING (.ZN (XNOR_1_4_N85_PULSESHAPING_OUT), .A1 (XNOR_1_3_N85_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_5_N85_PULSESHAPING (.ZN (XNOR_1_5_N85_PULSESHAPING_OUT), .A1 (XNOR_1_4_N85_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_6_N85_PULSESHAPING (.ZN (XNOR_1_6_N85_PULSESHAPING_OUT), .A1 (XNOR_1_5_N85_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_7_N85_PULSESHAPING (.ZN (N85), .A1 (XNOR_1_6_N85_PULSESHAPING_OUT), .A2 (GND));

      wire XNOR_1_1_N92_PULSESHAPING_OUT, XNOR_1_2_N92_PULSESHAPING_OUT, XNOR_1_3_N92_PULSESHAPING_OUT, XNOR_1_4_N92_PULSESHAPING_OUT, XNOR_1_5_N92_PULSESHAPING_OUT, XNOR_1_6_N92_PULSESHAPING_OUT;
      NOR2_X1 XNOR_1_1_N92_PULSESHAPING (.ZN (XNOR_1_1_N92_PULSESHAPING_OUT), .A1 (N92_PWL), .A2 (GND));
      NOR2_X1 XNOR_1_2_N92_PULSESHAPING (.ZN (XNOR_1_2_N92_PULSESHAPING_OUT), .A1 (XNOR_1_1_N92_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_3_N92_PULSESHAPING (.ZN (XNOR_1_3_N92_PULSESHAPING_OUT), .A1 (XNOR_1_2_N92_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_4_N92_PULSESHAPING (.ZN (XNOR_1_4_N92_PULSESHAPING_OUT), .A1 (XNOR_1_3_N92_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_5_N92_PULSESHAPING (.ZN (XNOR_1_5_N92_PULSESHAPING_OUT), .A1 (XNOR_1_4_N92_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_6_N92_PULSESHAPING (.ZN (XNOR_1_6_N92_PULSESHAPING_OUT), .A1 (XNOR_1_5_N92_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_7_N92_PULSESHAPING (.ZN (N92), .A1 (XNOR_1_6_N92_PULSESHAPING_OUT), .A2 (GND));

      wire XNOR_1_1_N99_PULSESHAPING_OUT, XNOR_1_2_N99_PULSESHAPING_OUT, XNOR_1_3_N99_PULSESHAPING_OUT, XNOR_1_4_N99_PULSESHAPING_OUT, XNOR_1_5_N99_PULSESHAPING_OUT, XNOR_1_6_N99_PULSESHAPING_OUT;
      NOR2_X1 XNOR_1_1_N99_PULSESHAPING (.ZN (XNOR_1_1_N99_PULSESHAPING_OUT), .A1 (N99_PWL), .A2 (GND));
      NOR2_X1 XNOR_1_2_N99_PULSESHAPING (.ZN (XNOR_1_2_N99_PULSESHAPING_OUT), .A1 (XNOR_1_1_N99_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_3_N99_PULSESHAPING (.ZN (XNOR_1_3_N99_PULSESHAPING_OUT), .A1 (XNOR_1_2_N99_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_4_N99_PULSESHAPING (.ZN (XNOR_1_4_N99_PULSESHAPING_OUT), .A1 (XNOR_1_3_N99_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_5_N99_PULSESHAPING (.ZN (XNOR_1_5_N99_PULSESHAPING_OUT), .A1 (XNOR_1_4_N99_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_6_N99_PULSESHAPING (.ZN (XNOR_1_6_N99_PULSESHAPING_OUT), .A1 (XNOR_1_5_N99_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_7_N99_PULSESHAPING (.ZN (N99), .A1 (XNOR_1_6_N99_PULSESHAPING_OUT), .A2 (GND));

      wire XNOR_1_1_N106_PULSESHAPING_OUT, XNOR_1_2_N106_PULSESHAPING_OUT, XNOR_1_3_N106_PULSESHAPING_OUT, XNOR_1_4_N106_PULSESHAPING_OUT, XNOR_1_5_N106_PULSESHAPING_OUT, XNOR_1_6_N106_PULSESHAPING_OUT;
      NOR2_X1 XNOR_1_1_N106_PULSESHAPING (.ZN (XNOR_1_1_N106_PULSESHAPING_OUT), .A1 (N106_PWL), .A2 (GND));
      NOR2_X1 XNOR_1_2_N106_PULSESHAPING (.ZN (XNOR_1_2_N106_PULSESHAPING_OUT), .A1 (XNOR_1_1_N106_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_3_N106_PULSESHAPING (.ZN (XNOR_1_3_N106_PULSESHAPING_OUT), .A1 (XNOR_1_2_N106_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_4_N106_PULSESHAPING (.ZN (XNOR_1_4_N106_PULSESHAPING_OUT), .A1 (XNOR_1_3_N106_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_5_N106_PULSESHAPING (.ZN (XNOR_1_5_N106_PULSESHAPING_OUT), .A1 (XNOR_1_4_N106_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_6_N106_PULSESHAPING (.ZN (XNOR_1_6_N106_PULSESHAPING_OUT), .A1 (XNOR_1_5_N106_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_7_N106_PULSESHAPING (.ZN (N106), .A1 (XNOR_1_6_N106_PULSESHAPING_OUT), .A2 (GND));

      wire XNOR_1_1_N113_PULSESHAPING_OUT, XNOR_1_2_N113_PULSESHAPING_OUT, XNOR_1_3_N113_PULSESHAPING_OUT, XNOR_1_4_N113_PULSESHAPING_OUT, XNOR_1_5_N113_PULSESHAPING_OUT, XNOR_1_6_N113_PULSESHAPING_OUT;
      NOR2_X1 XNOR_1_1_N113_PULSESHAPING (.ZN (XNOR_1_1_N113_PULSESHAPING_OUT), .A1 (N113_PWL), .A2 (GND));
      NOR2_X1 XNOR_1_2_N113_PULSESHAPING (.ZN (XNOR_1_2_N113_PULSESHAPING_OUT), .A1 (XNOR_1_1_N113_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_3_N113_PULSESHAPING (.ZN (XNOR_1_3_N113_PULSESHAPING_OUT), .A1 (XNOR_1_2_N113_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_4_N113_PULSESHAPING (.ZN (XNOR_1_4_N113_PULSESHAPING_OUT), .A1 (XNOR_1_3_N113_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_5_N113_PULSESHAPING (.ZN (XNOR_1_5_N113_PULSESHAPING_OUT), .A1 (XNOR_1_4_N113_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_6_N113_PULSESHAPING (.ZN (XNOR_1_6_N113_PULSESHAPING_OUT), .A1 (XNOR_1_5_N113_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_7_N113_PULSESHAPING (.ZN (N113), .A1 (XNOR_1_6_N113_PULSESHAPING_OUT), .A2 (GND));

      wire XNOR_1_1_N120_PULSESHAPING_OUT, XNOR_1_2_N120_PULSESHAPING_OUT, XNOR_1_3_N120_PULSESHAPING_OUT, XNOR_1_4_N120_PULSESHAPING_OUT, XNOR_1_5_N120_PULSESHAPING_OUT, XNOR_1_6_N120_PULSESHAPING_OUT;
      NOR2_X1 XNOR_1_1_N120_PULSESHAPING (.ZN (XNOR_1_1_N120_PULSESHAPING_OUT), .A1 (N120_PWL), .A2 (GND));
      NOR2_X1 XNOR_1_2_N120_PULSESHAPING (.ZN (XNOR_1_2_N120_PULSESHAPING_OUT), .A1 (XNOR_1_1_N120_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_3_N120_PULSESHAPING (.ZN (XNOR_1_3_N120_PULSESHAPING_OUT), .A1 (XNOR_1_2_N120_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_4_N120_PULSESHAPING (.ZN (XNOR_1_4_N120_PULSESHAPING_OUT), .A1 (XNOR_1_3_N120_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_5_N120_PULSESHAPING (.ZN (XNOR_1_5_N120_PULSESHAPING_OUT), .A1 (XNOR_1_4_N120_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_6_N120_PULSESHAPING (.ZN (XNOR_1_6_N120_PULSESHAPING_OUT), .A1 (XNOR_1_5_N120_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_7_N120_PULSESHAPING (.ZN (N120), .A1 (XNOR_1_6_N120_PULSESHAPING_OUT), .A2 (GND));

      wire XNOR_1_1_N127_PULSESHAPING_OUT, XNOR_1_2_N127_PULSESHAPING_OUT, XNOR_1_3_N127_PULSESHAPING_OUT, XNOR_1_4_N127_PULSESHAPING_OUT, XNOR_1_5_N127_PULSESHAPING_OUT, XNOR_1_6_N127_PULSESHAPING_OUT;
      NOR2_X1 XNOR_1_1_N127_PULSESHAPING (.ZN (XNOR_1_1_N127_PULSESHAPING_OUT), .A1 (N127_PWL), .A2 (GND));
      NOR2_X1 XNOR_1_2_N127_PULSESHAPING (.ZN (XNOR_1_2_N127_PULSESHAPING_OUT), .A1 (XNOR_1_1_N127_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_3_N127_PULSESHAPING (.ZN (XNOR_1_3_N127_PULSESHAPING_OUT), .A1 (XNOR_1_2_N127_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_4_N127_PULSESHAPING (.ZN (XNOR_1_4_N127_PULSESHAPING_OUT), .A1 (XNOR_1_3_N127_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_5_N127_PULSESHAPING (.ZN (XNOR_1_5_N127_PULSESHAPING_OUT), .A1 (XNOR_1_4_N127_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_6_N127_PULSESHAPING (.ZN (XNOR_1_6_N127_PULSESHAPING_OUT), .A1 (XNOR_1_5_N127_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_7_N127_PULSESHAPING (.ZN (N127), .A1 (XNOR_1_6_N127_PULSESHAPING_OUT), .A2 (GND));

      wire XNOR_1_1_N134_PULSESHAPING_OUT, XNOR_1_2_N134_PULSESHAPING_OUT, XNOR_1_3_N134_PULSESHAPING_OUT, XNOR_1_4_N134_PULSESHAPING_OUT, XNOR_1_5_N134_PULSESHAPING_OUT, XNOR_1_6_N134_PULSESHAPING_OUT;
      NOR2_X1 XNOR_1_1_N134_PULSESHAPING (.ZN (XNOR_1_1_N134_PULSESHAPING_OUT), .A1 (N134_PWL), .A2 (GND));
      NOR2_X1 XNOR_1_2_N134_PULSESHAPING (.ZN (XNOR_1_2_N134_PULSESHAPING_OUT), .A1 (XNOR_1_1_N134_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_3_N134_PULSESHAPING (.ZN (XNOR_1_3_N134_PULSESHAPING_OUT), .A1 (XNOR_1_2_N134_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_4_N134_PULSESHAPING (.ZN (XNOR_1_4_N134_PULSESHAPING_OUT), .A1 (XNOR_1_3_N134_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_5_N134_PULSESHAPING (.ZN (XNOR_1_5_N134_PULSESHAPING_OUT), .A1 (XNOR_1_4_N134_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_6_N134_PULSESHAPING (.ZN (XNOR_1_6_N134_PULSESHAPING_OUT), .A1 (XNOR_1_5_N134_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_7_N134_PULSESHAPING (.ZN (N134), .A1 (XNOR_1_6_N134_PULSESHAPING_OUT), .A2 (GND));

      wire XNOR_1_1_N141_PULSESHAPING_OUT, XNOR_1_2_N141_PULSESHAPING_OUT, XNOR_1_3_N141_PULSESHAPING_OUT, XNOR_1_4_N141_PULSESHAPING_OUT, XNOR_1_5_N141_PULSESHAPING_OUT, XNOR_1_6_N141_PULSESHAPING_OUT;
      NOR2_X1 XNOR_1_1_N141_PULSESHAPING (.ZN (XNOR_1_1_N141_PULSESHAPING_OUT), .A1 (N141_PWL), .A2 (GND));
      NOR2_X1 XNOR_1_2_N141_PULSESHAPING (.ZN (XNOR_1_2_N141_PULSESHAPING_OUT), .A1 (XNOR_1_1_N141_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_3_N141_PULSESHAPING (.ZN (XNOR_1_3_N141_PULSESHAPING_OUT), .A1 (XNOR_1_2_N141_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_4_N141_PULSESHAPING (.ZN (XNOR_1_4_N141_PULSESHAPING_OUT), .A1 (XNOR_1_3_N141_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_5_N141_PULSESHAPING (.ZN (XNOR_1_5_N141_PULSESHAPING_OUT), .A1 (XNOR_1_4_N141_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_6_N141_PULSESHAPING (.ZN (XNOR_1_6_N141_PULSESHAPING_OUT), .A1 (XNOR_1_5_N141_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_7_N141_PULSESHAPING (.ZN (N141), .A1 (XNOR_1_6_N141_PULSESHAPING_OUT), .A2 (GND));

      wire XNOR_1_1_N148_PULSESHAPING_OUT, XNOR_1_2_N148_PULSESHAPING_OUT, XNOR_1_3_N148_PULSESHAPING_OUT, XNOR_1_4_N148_PULSESHAPING_OUT, XNOR_1_5_N148_PULSESHAPING_OUT, XNOR_1_6_N148_PULSESHAPING_OUT;
      NOR2_X1 XNOR_1_1_N148_PULSESHAPING (.ZN (XNOR_1_1_N148_PULSESHAPING_OUT), .A1 (N148_PWL), .A2 (GND));
      NOR2_X1 XNOR_1_2_N148_PULSESHAPING (.ZN (XNOR_1_2_N148_PULSESHAPING_OUT), .A1 (XNOR_1_1_N148_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_3_N148_PULSESHAPING (.ZN (XNOR_1_3_N148_PULSESHAPING_OUT), .A1 (XNOR_1_2_N148_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_4_N148_PULSESHAPING (.ZN (XNOR_1_4_N148_PULSESHAPING_OUT), .A1 (XNOR_1_3_N148_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_5_N148_PULSESHAPING (.ZN (XNOR_1_5_N148_PULSESHAPING_OUT), .A1 (XNOR_1_4_N148_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_6_N148_PULSESHAPING (.ZN (XNOR_1_6_N148_PULSESHAPING_OUT), .A1 (XNOR_1_5_N148_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_7_N148_PULSESHAPING (.ZN (N148), .A1 (XNOR_1_6_N148_PULSESHAPING_OUT), .A2 (GND));

      wire XNOR_1_1_N155_PULSESHAPING_OUT, XNOR_1_2_N155_PULSESHAPING_OUT, XNOR_1_3_N155_PULSESHAPING_OUT, XNOR_1_4_N155_PULSESHAPING_OUT, XNOR_1_5_N155_PULSESHAPING_OUT, XNOR_1_6_N155_PULSESHAPING_OUT;
      NOR2_X1 XNOR_1_1_N155_PULSESHAPING (.ZN (XNOR_1_1_N155_PULSESHAPING_OUT), .A1 (N155_PWL), .A2 (GND));
      NOR2_X1 XNOR_1_2_N155_PULSESHAPING (.ZN (XNOR_1_2_N155_PULSESHAPING_OUT), .A1 (XNOR_1_1_N155_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_3_N155_PULSESHAPING (.ZN (XNOR_1_3_N155_PULSESHAPING_OUT), .A1 (XNOR_1_2_N155_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_4_N155_PULSESHAPING (.ZN (XNOR_1_4_N155_PULSESHAPING_OUT), .A1 (XNOR_1_3_N155_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_5_N155_PULSESHAPING (.ZN (XNOR_1_5_N155_PULSESHAPING_OUT), .A1 (XNOR_1_4_N155_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_6_N155_PULSESHAPING (.ZN (XNOR_1_6_N155_PULSESHAPING_OUT), .A1 (XNOR_1_5_N155_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_7_N155_PULSESHAPING (.ZN (N155), .A1 (XNOR_1_6_N155_PULSESHAPING_OUT), .A2 (GND));

      wire XNOR_1_1_N162_PULSESHAPING_OUT, XNOR_1_2_N162_PULSESHAPING_OUT, XNOR_1_3_N162_PULSESHAPING_OUT, XNOR_1_4_N162_PULSESHAPING_OUT, XNOR_1_5_N162_PULSESHAPING_OUT, XNOR_1_6_N162_PULSESHAPING_OUT;
      NOR2_X1 XNOR_1_1_N162_PULSESHAPING (.ZN (XNOR_1_1_N162_PULSESHAPING_OUT), .A1 (N162_PWL), .A2 (GND));
      NOR2_X1 XNOR_1_2_N162_PULSESHAPING (.ZN (XNOR_1_2_N162_PULSESHAPING_OUT), .A1 (XNOR_1_1_N162_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_3_N162_PULSESHAPING (.ZN (XNOR_1_3_N162_PULSESHAPING_OUT), .A1 (XNOR_1_2_N162_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_4_N162_PULSESHAPING (.ZN (XNOR_1_4_N162_PULSESHAPING_OUT), .A1 (XNOR_1_3_N162_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_5_N162_PULSESHAPING (.ZN (XNOR_1_5_N162_PULSESHAPING_OUT), .A1 (XNOR_1_4_N162_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_6_N162_PULSESHAPING (.ZN (XNOR_1_6_N162_PULSESHAPING_OUT), .A1 (XNOR_1_5_N162_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_7_N162_PULSESHAPING (.ZN (N162), .A1 (XNOR_1_6_N162_PULSESHAPING_OUT), .A2 (GND));

      wire XNOR_1_1_N169_PULSESHAPING_OUT, XNOR_1_2_N169_PULSESHAPING_OUT, XNOR_1_3_N169_PULSESHAPING_OUT, XNOR_1_4_N169_PULSESHAPING_OUT, XNOR_1_5_N169_PULSESHAPING_OUT, XNOR_1_6_N169_PULSESHAPING_OUT;
      NOR2_X1 XNOR_1_1_N169_PULSESHAPING (.ZN (XNOR_1_1_N169_PULSESHAPING_OUT), .A1 (N169_PWL), .A2 (GND));
      NOR2_X1 XNOR_1_2_N169_PULSESHAPING (.ZN (XNOR_1_2_N169_PULSESHAPING_OUT), .A1 (XNOR_1_1_N169_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_3_N169_PULSESHAPING (.ZN (XNOR_1_3_N169_PULSESHAPING_OUT), .A1 (XNOR_1_2_N169_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_4_N169_PULSESHAPING (.ZN (XNOR_1_4_N169_PULSESHAPING_OUT), .A1 (XNOR_1_3_N169_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_5_N169_PULSESHAPING (.ZN (XNOR_1_5_N169_PULSESHAPING_OUT), .A1 (XNOR_1_4_N169_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_6_N169_PULSESHAPING (.ZN (XNOR_1_6_N169_PULSESHAPING_OUT), .A1 (XNOR_1_5_N169_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_7_N169_PULSESHAPING (.ZN (N169), .A1 (XNOR_1_6_N169_PULSESHAPING_OUT), .A2 (GND));

      wire XNOR_1_1_N176_PULSESHAPING_OUT, XNOR_1_2_N176_PULSESHAPING_OUT, XNOR_1_3_N176_PULSESHAPING_OUT, XNOR_1_4_N176_PULSESHAPING_OUT, XNOR_1_5_N176_PULSESHAPING_OUT, XNOR_1_6_N176_PULSESHAPING_OUT;
      NOR2_X1 XNOR_1_1_N176_PULSESHAPING (.ZN (XNOR_1_1_N176_PULSESHAPING_OUT), .A1 (N176_PWL), .A2 (GND));
      NOR2_X1 XNOR_1_2_N176_PULSESHAPING (.ZN (XNOR_1_2_N176_PULSESHAPING_OUT), .A1 (XNOR_1_1_N176_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_3_N176_PULSESHAPING (.ZN (XNOR_1_3_N176_PULSESHAPING_OUT), .A1 (XNOR_1_2_N176_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_4_N176_PULSESHAPING (.ZN (XNOR_1_4_N176_PULSESHAPING_OUT), .A1 (XNOR_1_3_N176_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_5_N176_PULSESHAPING (.ZN (XNOR_1_5_N176_PULSESHAPING_OUT), .A1 (XNOR_1_4_N176_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_6_N176_PULSESHAPING (.ZN (XNOR_1_6_N176_PULSESHAPING_OUT), .A1 (XNOR_1_5_N176_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_7_N176_PULSESHAPING (.ZN (N176), .A1 (XNOR_1_6_N176_PULSESHAPING_OUT), .A2 (GND));

      wire XNOR_1_1_N183_PULSESHAPING_OUT, XNOR_1_2_N183_PULSESHAPING_OUT, XNOR_1_3_N183_PULSESHAPING_OUT, XNOR_1_4_N183_PULSESHAPING_OUT, XNOR_1_5_N183_PULSESHAPING_OUT, XNOR_1_6_N183_PULSESHAPING_OUT;
      NOR2_X1 XNOR_1_1_N183_PULSESHAPING (.ZN (XNOR_1_1_N183_PULSESHAPING_OUT), .A1 (N183_PWL), .A2 (GND));
      NOR2_X1 XNOR_1_2_N183_PULSESHAPING (.ZN (XNOR_1_2_N183_PULSESHAPING_OUT), .A1 (XNOR_1_1_N183_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_3_N183_PULSESHAPING (.ZN (XNOR_1_3_N183_PULSESHAPING_OUT), .A1 (XNOR_1_2_N183_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_4_N183_PULSESHAPING (.ZN (XNOR_1_4_N183_PULSESHAPING_OUT), .A1 (XNOR_1_3_N183_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_5_N183_PULSESHAPING (.ZN (XNOR_1_5_N183_PULSESHAPING_OUT), .A1 (XNOR_1_4_N183_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_6_N183_PULSESHAPING (.ZN (XNOR_1_6_N183_PULSESHAPING_OUT), .A1 (XNOR_1_5_N183_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_7_N183_PULSESHAPING (.ZN (N183), .A1 (XNOR_1_6_N183_PULSESHAPING_OUT), .A2 (GND));

      wire XNOR_1_1_N190_PULSESHAPING_OUT, XNOR_1_2_N190_PULSESHAPING_OUT, XNOR_1_3_N190_PULSESHAPING_OUT, XNOR_1_4_N190_PULSESHAPING_OUT, XNOR_1_5_N190_PULSESHAPING_OUT, XNOR_1_6_N190_PULSESHAPING_OUT;
      NOR2_X1 XNOR_1_1_N190_PULSESHAPING (.ZN (XNOR_1_1_N190_PULSESHAPING_OUT), .A1 (N190_PWL), .A2 (GND));
      NOR2_X1 XNOR_1_2_N190_PULSESHAPING (.ZN (XNOR_1_2_N190_PULSESHAPING_OUT), .A1 (XNOR_1_1_N190_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_3_N190_PULSESHAPING (.ZN (XNOR_1_3_N190_PULSESHAPING_OUT), .A1 (XNOR_1_2_N190_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_4_N190_PULSESHAPING (.ZN (XNOR_1_4_N190_PULSESHAPING_OUT), .A1 (XNOR_1_3_N190_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_5_N190_PULSESHAPING (.ZN (XNOR_1_5_N190_PULSESHAPING_OUT), .A1 (XNOR_1_4_N190_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_6_N190_PULSESHAPING (.ZN (XNOR_1_6_N190_PULSESHAPING_OUT), .A1 (XNOR_1_5_N190_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_7_N190_PULSESHAPING (.ZN (N190), .A1 (XNOR_1_6_N190_PULSESHAPING_OUT), .A2 (GND));

      wire XNOR_1_1_N197_PULSESHAPING_OUT, XNOR_1_2_N197_PULSESHAPING_OUT, XNOR_1_3_N197_PULSESHAPING_OUT, XNOR_1_4_N197_PULSESHAPING_OUT, XNOR_1_5_N197_PULSESHAPING_OUT, XNOR_1_6_N197_PULSESHAPING_OUT;
      NOR2_X1 XNOR_1_1_N197_PULSESHAPING (.ZN (XNOR_1_1_N197_PULSESHAPING_OUT), .A1 (N197_PWL), .A2 (GND));
      NOR2_X1 XNOR_1_2_N197_PULSESHAPING (.ZN (XNOR_1_2_N197_PULSESHAPING_OUT), .A1 (XNOR_1_1_N197_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_3_N197_PULSESHAPING (.ZN (XNOR_1_3_N197_PULSESHAPING_OUT), .A1 (XNOR_1_2_N197_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_4_N197_PULSESHAPING (.ZN (XNOR_1_4_N197_PULSESHAPING_OUT), .A1 (XNOR_1_3_N197_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_5_N197_PULSESHAPING (.ZN (XNOR_1_5_N197_PULSESHAPING_OUT), .A1 (XNOR_1_4_N197_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_6_N197_PULSESHAPING (.ZN (XNOR_1_6_N197_PULSESHAPING_OUT), .A1 (XNOR_1_5_N197_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_7_N197_PULSESHAPING (.ZN (N197), .A1 (XNOR_1_6_N197_PULSESHAPING_OUT), .A2 (GND));

      wire XNOR_1_1_N204_PULSESHAPING_OUT, XNOR_1_2_N204_PULSESHAPING_OUT, XNOR_1_3_N204_PULSESHAPING_OUT, XNOR_1_4_N204_PULSESHAPING_OUT, XNOR_1_5_N204_PULSESHAPING_OUT, XNOR_1_6_N204_PULSESHAPING_OUT;
      NOR2_X1 XNOR_1_1_N204_PULSESHAPING (.ZN (XNOR_1_1_N204_PULSESHAPING_OUT), .A1 (N204_PWL), .A2 (GND));
      NOR2_X1 XNOR_1_2_N204_PULSESHAPING (.ZN (XNOR_1_2_N204_PULSESHAPING_OUT), .A1 (XNOR_1_1_N204_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_3_N204_PULSESHAPING (.ZN (XNOR_1_3_N204_PULSESHAPING_OUT), .A1 (XNOR_1_2_N204_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_4_N204_PULSESHAPING (.ZN (XNOR_1_4_N204_PULSESHAPING_OUT), .A1 (XNOR_1_3_N204_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_5_N204_PULSESHAPING (.ZN (XNOR_1_5_N204_PULSESHAPING_OUT), .A1 (XNOR_1_4_N204_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_6_N204_PULSESHAPING (.ZN (XNOR_1_6_N204_PULSESHAPING_OUT), .A1 (XNOR_1_5_N204_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_7_N204_PULSESHAPING (.ZN (N204), .A1 (XNOR_1_6_N204_PULSESHAPING_OUT), .A2 (GND));

      wire XNOR_1_1_N211_PULSESHAPING_OUT, XNOR_1_2_N211_PULSESHAPING_OUT, XNOR_1_3_N211_PULSESHAPING_OUT, XNOR_1_4_N211_PULSESHAPING_OUT, XNOR_1_5_N211_PULSESHAPING_OUT, XNOR_1_6_N211_PULSESHAPING_OUT;
      NOR2_X1 XNOR_1_1_N211_PULSESHAPING (.ZN (XNOR_1_1_N211_PULSESHAPING_OUT), .A1 (N211_PWL), .A2 (GND));
      NOR2_X1 XNOR_1_2_N211_PULSESHAPING (.ZN (XNOR_1_2_N211_PULSESHAPING_OUT), .A1 (XNOR_1_1_N211_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_3_N211_PULSESHAPING (.ZN (XNOR_1_3_N211_PULSESHAPING_OUT), .A1 (XNOR_1_2_N211_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_4_N211_PULSESHAPING (.ZN (XNOR_1_4_N211_PULSESHAPING_OUT), .A1 (XNOR_1_3_N211_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_5_N211_PULSESHAPING (.ZN (XNOR_1_5_N211_PULSESHAPING_OUT), .A1 (XNOR_1_4_N211_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_6_N211_PULSESHAPING (.ZN (XNOR_1_6_N211_PULSESHAPING_OUT), .A1 (XNOR_1_5_N211_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_7_N211_PULSESHAPING (.ZN (N211), .A1 (XNOR_1_6_N211_PULSESHAPING_OUT), .A2 (GND));

      wire XNOR_1_1_N218_PULSESHAPING_OUT, XNOR_1_2_N218_PULSESHAPING_OUT, XNOR_1_3_N218_PULSESHAPING_OUT, XNOR_1_4_N218_PULSESHAPING_OUT, XNOR_1_5_N218_PULSESHAPING_OUT, XNOR_1_6_N218_PULSESHAPING_OUT;
      NOR2_X1 XNOR_1_1_N218_PULSESHAPING (.ZN (XNOR_1_1_N218_PULSESHAPING_OUT), .A1 (N218_PWL), .A2 (GND));
      NOR2_X1 XNOR_1_2_N218_PULSESHAPING (.ZN (XNOR_1_2_N218_PULSESHAPING_OUT), .A1 (XNOR_1_1_N218_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_3_N218_PULSESHAPING (.ZN (XNOR_1_3_N218_PULSESHAPING_OUT), .A1 (XNOR_1_2_N218_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_4_N218_PULSESHAPING (.ZN (XNOR_1_4_N218_PULSESHAPING_OUT), .A1 (XNOR_1_3_N218_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_5_N218_PULSESHAPING (.ZN (XNOR_1_5_N218_PULSESHAPING_OUT), .A1 (XNOR_1_4_N218_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_6_N218_PULSESHAPING (.ZN (XNOR_1_6_N218_PULSESHAPING_OUT), .A1 (XNOR_1_5_N218_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_7_N218_PULSESHAPING (.ZN (N218), .A1 (XNOR_1_6_N218_PULSESHAPING_OUT), .A2 (GND));

      wire XNOR_1_1_N225_PULSESHAPING_OUT, XNOR_1_2_N225_PULSESHAPING_OUT, XNOR_1_3_N225_PULSESHAPING_OUT, XNOR_1_4_N225_PULSESHAPING_OUT, XNOR_1_5_N225_PULSESHAPING_OUT, XNOR_1_6_N225_PULSESHAPING_OUT;
      NOR2_X1 XNOR_1_1_N225_PULSESHAPING (.ZN (XNOR_1_1_N225_PULSESHAPING_OUT), .A1 (N225_PWL), .A2 (GND));
      NOR2_X1 XNOR_1_2_N225_PULSESHAPING (.ZN (XNOR_1_2_N225_PULSESHAPING_OUT), .A1 (XNOR_1_1_N225_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_3_N225_PULSESHAPING (.ZN (XNOR_1_3_N225_PULSESHAPING_OUT), .A1 (XNOR_1_2_N225_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_4_N225_PULSESHAPING (.ZN (XNOR_1_4_N225_PULSESHAPING_OUT), .A1 (XNOR_1_3_N225_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_5_N225_PULSESHAPING (.ZN (XNOR_1_5_N225_PULSESHAPING_OUT), .A1 (XNOR_1_4_N225_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_6_N225_PULSESHAPING (.ZN (XNOR_1_6_N225_PULSESHAPING_OUT), .A1 (XNOR_1_5_N225_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_7_N225_PULSESHAPING (.ZN (N225), .A1 (XNOR_1_6_N225_PULSESHAPING_OUT), .A2 (GND));

      wire XNOR_1_1_N226_PULSESHAPING_OUT, XNOR_1_2_N226_PULSESHAPING_OUT, XNOR_1_3_N226_PULSESHAPING_OUT, XNOR_1_4_N226_PULSESHAPING_OUT, XNOR_1_5_N226_PULSESHAPING_OUT, XNOR_1_6_N226_PULSESHAPING_OUT;
      NOR2_X1 XNOR_1_1_N226_PULSESHAPING (.ZN (XNOR_1_1_N226_PULSESHAPING_OUT), .A1 (N226_PWL), .A2 (GND));
      NOR2_X1 XNOR_1_2_N226_PULSESHAPING (.ZN (XNOR_1_2_N226_PULSESHAPING_OUT), .A1 (XNOR_1_1_N226_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_3_N226_PULSESHAPING (.ZN (XNOR_1_3_N226_PULSESHAPING_OUT), .A1 (XNOR_1_2_N226_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_4_N226_PULSESHAPING (.ZN (XNOR_1_4_N226_PULSESHAPING_OUT), .A1 (XNOR_1_3_N226_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_5_N226_PULSESHAPING (.ZN (XNOR_1_5_N226_PULSESHAPING_OUT), .A1 (XNOR_1_4_N226_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_6_N226_PULSESHAPING (.ZN (XNOR_1_6_N226_PULSESHAPING_OUT), .A1 (XNOR_1_5_N226_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_7_N226_PULSESHAPING (.ZN (N226), .A1 (XNOR_1_6_N226_PULSESHAPING_OUT), .A2 (GND));

      wire XNOR_1_1_N227_PULSESHAPING_OUT, XNOR_1_2_N227_PULSESHAPING_OUT, XNOR_1_3_N227_PULSESHAPING_OUT, XNOR_1_4_N227_PULSESHAPING_OUT, XNOR_1_5_N227_PULSESHAPING_OUT, XNOR_1_6_N227_PULSESHAPING_OUT;
      NOR2_X1 XNOR_1_1_N227_PULSESHAPING (.ZN (XNOR_1_1_N227_PULSESHAPING_OUT), .A1 (N227_PWL), .A2 (GND));
      NOR2_X1 XNOR_1_2_N227_PULSESHAPING (.ZN (XNOR_1_2_N227_PULSESHAPING_OUT), .A1 (XNOR_1_1_N227_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_3_N227_PULSESHAPING (.ZN (XNOR_1_3_N227_PULSESHAPING_OUT), .A1 (XNOR_1_2_N227_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_4_N227_PULSESHAPING (.ZN (XNOR_1_4_N227_PULSESHAPING_OUT), .A1 (XNOR_1_3_N227_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_5_N227_PULSESHAPING (.ZN (XNOR_1_5_N227_PULSESHAPING_OUT), .A1 (XNOR_1_4_N227_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_6_N227_PULSESHAPING (.ZN (XNOR_1_6_N227_PULSESHAPING_OUT), .A1 (XNOR_1_5_N227_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_7_N227_PULSESHAPING (.ZN (N227), .A1 (XNOR_1_6_N227_PULSESHAPING_OUT), .A2 (GND));

      wire XNOR_1_1_N228_PULSESHAPING_OUT, XNOR_1_2_N228_PULSESHAPING_OUT, XNOR_1_3_N228_PULSESHAPING_OUT, XNOR_1_4_N228_PULSESHAPING_OUT, XNOR_1_5_N228_PULSESHAPING_OUT, XNOR_1_6_N228_PULSESHAPING_OUT;
      NOR2_X1 XNOR_1_1_N228_PULSESHAPING (.ZN (XNOR_1_1_N228_PULSESHAPING_OUT), .A1 (N228_PWL), .A2 (GND));
      NOR2_X1 XNOR_1_2_N228_PULSESHAPING (.ZN (XNOR_1_2_N228_PULSESHAPING_OUT), .A1 (XNOR_1_1_N228_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_3_N228_PULSESHAPING (.ZN (XNOR_1_3_N228_PULSESHAPING_OUT), .A1 (XNOR_1_2_N228_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_4_N228_PULSESHAPING (.ZN (XNOR_1_4_N228_PULSESHAPING_OUT), .A1 (XNOR_1_3_N228_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_5_N228_PULSESHAPING (.ZN (XNOR_1_5_N228_PULSESHAPING_OUT), .A1 (XNOR_1_4_N228_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_6_N228_PULSESHAPING (.ZN (XNOR_1_6_N228_PULSESHAPING_OUT), .A1 (XNOR_1_5_N228_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_7_N228_PULSESHAPING (.ZN (N228), .A1 (XNOR_1_6_N228_PULSESHAPING_OUT), .A2 (GND));

      wire XNOR_1_1_N229_PULSESHAPING_OUT, XNOR_1_2_N229_PULSESHAPING_OUT, XNOR_1_3_N229_PULSESHAPING_OUT, XNOR_1_4_N229_PULSESHAPING_OUT, XNOR_1_5_N229_PULSESHAPING_OUT, XNOR_1_6_N229_PULSESHAPING_OUT;
      NOR2_X1 XNOR_1_1_N229_PULSESHAPING (.ZN (XNOR_1_1_N229_PULSESHAPING_OUT), .A1 (N229_PWL), .A2 (GND));
      NOR2_X1 XNOR_1_2_N229_PULSESHAPING (.ZN (XNOR_1_2_N229_PULSESHAPING_OUT), .A1 (XNOR_1_1_N229_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_3_N229_PULSESHAPING (.ZN (XNOR_1_3_N229_PULSESHAPING_OUT), .A1 (XNOR_1_2_N229_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_4_N229_PULSESHAPING (.ZN (XNOR_1_4_N229_PULSESHAPING_OUT), .A1 (XNOR_1_3_N229_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_5_N229_PULSESHAPING (.ZN (XNOR_1_5_N229_PULSESHAPING_OUT), .A1 (XNOR_1_4_N229_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_6_N229_PULSESHAPING (.ZN (XNOR_1_6_N229_PULSESHAPING_OUT), .A1 (XNOR_1_5_N229_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_7_N229_PULSESHAPING (.ZN (N229), .A1 (XNOR_1_6_N229_PULSESHAPING_OUT), .A2 (GND));

      wire XNOR_1_1_N230_PULSESHAPING_OUT, XNOR_1_2_N230_PULSESHAPING_OUT, XNOR_1_3_N230_PULSESHAPING_OUT, XNOR_1_4_N230_PULSESHAPING_OUT, XNOR_1_5_N230_PULSESHAPING_OUT, XNOR_1_6_N230_PULSESHAPING_OUT;
      NOR2_X1 XNOR_1_1_N230_PULSESHAPING (.ZN (XNOR_1_1_N230_PULSESHAPING_OUT), .A1 (N230_PWL), .A2 (GND));
      NOR2_X1 XNOR_1_2_N230_PULSESHAPING (.ZN (XNOR_1_2_N230_PULSESHAPING_OUT), .A1 (XNOR_1_1_N230_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_3_N230_PULSESHAPING (.ZN (XNOR_1_3_N230_PULSESHAPING_OUT), .A1 (XNOR_1_2_N230_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_4_N230_PULSESHAPING (.ZN (XNOR_1_4_N230_PULSESHAPING_OUT), .A1 (XNOR_1_3_N230_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_5_N230_PULSESHAPING (.ZN (XNOR_1_5_N230_PULSESHAPING_OUT), .A1 (XNOR_1_4_N230_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_6_N230_PULSESHAPING (.ZN (XNOR_1_6_N230_PULSESHAPING_OUT), .A1 (XNOR_1_5_N230_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_7_N230_PULSESHAPING (.ZN (N230), .A1 (XNOR_1_6_N230_PULSESHAPING_OUT), .A2 (GND));

      wire XNOR_1_1_N231_PULSESHAPING_OUT, XNOR_1_2_N231_PULSESHAPING_OUT, XNOR_1_3_N231_PULSESHAPING_OUT, XNOR_1_4_N231_PULSESHAPING_OUT, XNOR_1_5_N231_PULSESHAPING_OUT, XNOR_1_6_N231_PULSESHAPING_OUT;
      NOR2_X1 XNOR_1_1_N231_PULSESHAPING (.ZN (XNOR_1_1_N231_PULSESHAPING_OUT), .A1 (N231_PWL), .A2 (GND));
      NOR2_X1 XNOR_1_2_N231_PULSESHAPING (.ZN (XNOR_1_2_N231_PULSESHAPING_OUT), .A1 (XNOR_1_1_N231_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_3_N231_PULSESHAPING (.ZN (XNOR_1_3_N231_PULSESHAPING_OUT), .A1 (XNOR_1_2_N231_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_4_N231_PULSESHAPING (.ZN (XNOR_1_4_N231_PULSESHAPING_OUT), .A1 (XNOR_1_3_N231_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_5_N231_PULSESHAPING (.ZN (XNOR_1_5_N231_PULSESHAPING_OUT), .A1 (XNOR_1_4_N231_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_6_N231_PULSESHAPING (.ZN (XNOR_1_6_N231_PULSESHAPING_OUT), .A1 (XNOR_1_5_N231_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_7_N231_PULSESHAPING (.ZN (N231), .A1 (XNOR_1_6_N231_PULSESHAPING_OUT), .A2 (GND));

      wire XNOR_1_1_N232_PULSESHAPING_OUT, XNOR_1_2_N232_PULSESHAPING_OUT, XNOR_1_3_N232_PULSESHAPING_OUT, XNOR_1_4_N232_PULSESHAPING_OUT, XNOR_1_5_N232_PULSESHAPING_OUT, XNOR_1_6_N232_PULSESHAPING_OUT;
      NOR2_X1 XNOR_1_1_N232_PULSESHAPING (.ZN (XNOR_1_1_N232_PULSESHAPING_OUT), .A1 (N232_PWL), .A2 (GND));
      NOR2_X1 XNOR_1_2_N232_PULSESHAPING (.ZN (XNOR_1_2_N232_PULSESHAPING_OUT), .A1 (XNOR_1_1_N232_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_3_N232_PULSESHAPING (.ZN (XNOR_1_3_N232_PULSESHAPING_OUT), .A1 (XNOR_1_2_N232_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_4_N232_PULSESHAPING (.ZN (XNOR_1_4_N232_PULSESHAPING_OUT), .A1 (XNOR_1_3_N232_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_5_N232_PULSESHAPING (.ZN (XNOR_1_5_N232_PULSESHAPING_OUT), .A1 (XNOR_1_4_N232_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_6_N232_PULSESHAPING (.ZN (XNOR_1_6_N232_PULSESHAPING_OUT), .A1 (XNOR_1_5_N232_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_7_N232_PULSESHAPING (.ZN (N232), .A1 (XNOR_1_6_N232_PULSESHAPING_OUT), .A2 (GND));

      wire XNOR_1_1_N233_PULSESHAPING_OUT, XNOR_1_2_N233_PULSESHAPING_OUT, XNOR_1_3_N233_PULSESHAPING_OUT, XNOR_1_4_N233_PULSESHAPING_OUT, XNOR_1_5_N233_PULSESHAPING_OUT, XNOR_1_6_N233_PULSESHAPING_OUT;
      NOR2_X1 XNOR_1_1_N233_PULSESHAPING (.ZN (XNOR_1_1_N233_PULSESHAPING_OUT), .A1 (N233_PWL), .A2 (GND));
      NOR2_X1 XNOR_1_2_N233_PULSESHAPING (.ZN (XNOR_1_2_N233_PULSESHAPING_OUT), .A1 (XNOR_1_1_N233_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_3_N233_PULSESHAPING (.ZN (XNOR_1_3_N233_PULSESHAPING_OUT), .A1 (XNOR_1_2_N233_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_4_N233_PULSESHAPING (.ZN (XNOR_1_4_N233_PULSESHAPING_OUT), .A1 (XNOR_1_3_N233_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_5_N233_PULSESHAPING (.ZN (XNOR_1_5_N233_PULSESHAPING_OUT), .A1 (XNOR_1_4_N233_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_6_N233_PULSESHAPING (.ZN (XNOR_1_6_N233_PULSESHAPING_OUT), .A1 (XNOR_1_5_N233_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_7_N233_PULSESHAPING (.ZN (N233), .A1 (XNOR_1_6_N233_PULSESHAPING_OUT), .A2 (GND));



      wire XNOR_1_1_AND2_NUM0_OUT, XNOR_1_2_AND2_NUM0_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM0 (.ZN (XNOR_1_1_AND2_NUM0_OUT), .A1 (N225), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM0 (.ZN (XNOR_1_2_AND2_NUM0_OUT), .A1 (GND), .A2 (N233));
      NOR2_X1 XNOR_1_3_AND2_NUM0 (.ZN (N242), .A1 (XNOR_1_1_AND2_NUM0_OUT), .A2 (XNOR_1_2_AND2_NUM0_OUT));
      wire XNOR_1_1_AND2_NUM1_OUT, XNOR_1_2_AND2_NUM1_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM1 (.ZN (XNOR_1_1_AND2_NUM1_OUT), .A1 (N226), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM1 (.ZN (XNOR_1_2_AND2_NUM1_OUT), .A1 (GND), .A2 (N233));
      NOR2_X1 XNOR_1_3_AND2_NUM1 (.ZN (N245), .A1 (XNOR_1_1_AND2_NUM1_OUT), .A2 (XNOR_1_2_AND2_NUM1_OUT));
      wire XNOR_1_1_AND2_NUM2_OUT, XNOR_1_2_AND2_NUM2_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM2 (.ZN (XNOR_1_1_AND2_NUM2_OUT), .A1 (N227), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM2 (.ZN (XNOR_1_2_AND2_NUM2_OUT), .A1 (GND), .A2 (N233));
      NOR2_X1 XNOR_1_3_AND2_NUM2 (.ZN (N248), .A1 (XNOR_1_1_AND2_NUM2_OUT), .A2 (XNOR_1_2_AND2_NUM2_OUT));
      wire XNOR_1_1_AND2_NUM3_OUT, XNOR_1_2_AND2_NUM3_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM3 (.ZN (XNOR_1_1_AND2_NUM3_OUT), .A1 (N228), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM3 (.ZN (XNOR_1_2_AND2_NUM3_OUT), .A1 (GND), .A2 (N233));
      NOR2_X1 XNOR_1_3_AND2_NUM3 (.ZN (N251), .A1 (XNOR_1_1_AND2_NUM3_OUT), .A2 (XNOR_1_2_AND2_NUM3_OUT));
      wire XNOR_1_1_AND2_NUM4_OUT, XNOR_1_2_AND2_NUM4_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM4 (.ZN (XNOR_1_1_AND2_NUM4_OUT), .A1 (N229), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM4 (.ZN (XNOR_1_2_AND2_NUM4_OUT), .A1 (GND), .A2 (N233));
      NOR2_X1 XNOR_1_3_AND2_NUM4 (.ZN (N254), .A1 (XNOR_1_1_AND2_NUM4_OUT), .A2 (XNOR_1_2_AND2_NUM4_OUT));
      wire XNOR_1_1_AND2_NUM5_OUT, XNOR_1_2_AND2_NUM5_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM5 (.ZN (XNOR_1_1_AND2_NUM5_OUT), .A1 (N230), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM5 (.ZN (XNOR_1_2_AND2_NUM5_OUT), .A1 (GND), .A2 (N233));
      NOR2_X1 XNOR_1_3_AND2_NUM5 (.ZN (N257), .A1 (XNOR_1_1_AND2_NUM5_OUT), .A2 (XNOR_1_2_AND2_NUM5_OUT));
      wire XNOR_1_1_AND2_NUM6_OUT, XNOR_1_2_AND2_NUM6_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM6 (.ZN (XNOR_1_1_AND2_NUM6_OUT), .A1 (N231), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM6 (.ZN (XNOR_1_2_AND2_NUM6_OUT), .A1 (GND), .A2 (N233));
      NOR2_X1 XNOR_1_3_AND2_NUM6 (.ZN (N260), .A1 (XNOR_1_1_AND2_NUM6_OUT), .A2 (XNOR_1_2_AND2_NUM6_OUT));
      wire XNOR_1_1_AND2_NUM7_OUT, XNOR_1_2_AND2_NUM7_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM7 (.ZN (XNOR_1_1_AND2_NUM7_OUT), .A1 (N232), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM7 (.ZN (XNOR_1_2_AND2_NUM7_OUT), .A1 (GND), .A2 (N233));
      NOR2_X1 XNOR_1_3_AND2_NUM7 (.ZN (N263), .A1 (XNOR_1_1_AND2_NUM7_OUT), .A2 (XNOR_1_2_AND2_NUM7_OUT));
      wire XNOR_1_1_NAND2_NUM0_OUT, XNOR_1_2_NAND2_NUM0_OUT, XNOR_1_3_NAND2_NUM0_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM0 (.ZN (XNOR_1_1_NAND2_NUM0_OUT), .A1 (N1), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM0 (.ZN (XNOR_1_2_NAND2_NUM0_OUT), .A1 (GND), .A2 (N8));
      NOR2_X1 XNOR_1_3_NAND2_NUM0 (.ZN (XNOR_1_3_NAND2_NUM0_OUT), .A1 (XNOR_1_1_NAND2_NUM0_OUT), .A2 (XNOR_1_2_NAND2_NUM0_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM0 (.ZN (N266), .A1 (XNOR_1_3_NAND2_NUM0_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM1_OUT, XNOR_1_2_NAND2_NUM1_OUT, XNOR_1_3_NAND2_NUM1_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM1 (.ZN (XNOR_1_1_NAND2_NUM1_OUT), .A1 (N15), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM1 (.ZN (XNOR_1_2_NAND2_NUM1_OUT), .A1 (GND), .A2 (N22));
      NOR2_X1 XNOR_1_3_NAND2_NUM1 (.ZN (XNOR_1_3_NAND2_NUM1_OUT), .A1 (XNOR_1_1_NAND2_NUM1_OUT), .A2 (XNOR_1_2_NAND2_NUM1_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM1 (.ZN (N269), .A1 (XNOR_1_3_NAND2_NUM1_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM2_OUT, XNOR_1_2_NAND2_NUM2_OUT, XNOR_1_3_NAND2_NUM2_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM2 (.ZN (XNOR_1_1_NAND2_NUM2_OUT), .A1 (N29), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM2 (.ZN (XNOR_1_2_NAND2_NUM2_OUT), .A1 (GND), .A2 (N36));
      NOR2_X1 XNOR_1_3_NAND2_NUM2 (.ZN (XNOR_1_3_NAND2_NUM2_OUT), .A1 (XNOR_1_1_NAND2_NUM2_OUT), .A2 (XNOR_1_2_NAND2_NUM2_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM2 (.ZN (N272), .A1 (XNOR_1_3_NAND2_NUM2_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM3_OUT, XNOR_1_2_NAND2_NUM3_OUT, XNOR_1_3_NAND2_NUM3_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM3 (.ZN (XNOR_1_1_NAND2_NUM3_OUT), .A1 (N43), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM3 (.ZN (XNOR_1_2_NAND2_NUM3_OUT), .A1 (GND), .A2 (N50));
      NOR2_X1 XNOR_1_3_NAND2_NUM3 (.ZN (XNOR_1_3_NAND2_NUM3_OUT), .A1 (XNOR_1_1_NAND2_NUM3_OUT), .A2 (XNOR_1_2_NAND2_NUM3_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM3 (.ZN (N275), .A1 (XNOR_1_3_NAND2_NUM3_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM4_OUT, XNOR_1_2_NAND2_NUM4_OUT, XNOR_1_3_NAND2_NUM4_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM4 (.ZN (XNOR_1_1_NAND2_NUM4_OUT), .A1 (N57), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM4 (.ZN (XNOR_1_2_NAND2_NUM4_OUT), .A1 (GND), .A2 (N64));
      NOR2_X1 XNOR_1_3_NAND2_NUM4 (.ZN (XNOR_1_3_NAND2_NUM4_OUT), .A1 (XNOR_1_1_NAND2_NUM4_OUT), .A2 (XNOR_1_2_NAND2_NUM4_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM4 (.ZN (N278), .A1 (XNOR_1_3_NAND2_NUM4_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM5_OUT, XNOR_1_2_NAND2_NUM5_OUT, XNOR_1_3_NAND2_NUM5_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM5 (.ZN (XNOR_1_1_NAND2_NUM5_OUT), .A1 (N71), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM5 (.ZN (XNOR_1_2_NAND2_NUM5_OUT), .A1 (GND), .A2 (N78));
      NOR2_X1 XNOR_1_3_NAND2_NUM5 (.ZN (XNOR_1_3_NAND2_NUM5_OUT), .A1 (XNOR_1_1_NAND2_NUM5_OUT), .A2 (XNOR_1_2_NAND2_NUM5_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM5 (.ZN (N281), .A1 (XNOR_1_3_NAND2_NUM5_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM6_OUT, XNOR_1_2_NAND2_NUM6_OUT, XNOR_1_3_NAND2_NUM6_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM6 (.ZN (XNOR_1_1_NAND2_NUM6_OUT), .A1 (N85), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM6 (.ZN (XNOR_1_2_NAND2_NUM6_OUT), .A1 (GND), .A2 (N92));
      NOR2_X1 XNOR_1_3_NAND2_NUM6 (.ZN (XNOR_1_3_NAND2_NUM6_OUT), .A1 (XNOR_1_1_NAND2_NUM6_OUT), .A2 (XNOR_1_2_NAND2_NUM6_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM6 (.ZN (N284), .A1 (XNOR_1_3_NAND2_NUM6_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM7_OUT, XNOR_1_2_NAND2_NUM7_OUT, XNOR_1_3_NAND2_NUM7_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM7 (.ZN (XNOR_1_1_NAND2_NUM7_OUT), .A1 (N99), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM7 (.ZN (XNOR_1_2_NAND2_NUM7_OUT), .A1 (GND), .A2 (N106));
      NOR2_X1 XNOR_1_3_NAND2_NUM7 (.ZN (XNOR_1_3_NAND2_NUM7_OUT), .A1 (XNOR_1_1_NAND2_NUM7_OUT), .A2 (XNOR_1_2_NAND2_NUM7_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM7 (.ZN (N287), .A1 (XNOR_1_3_NAND2_NUM7_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM8_OUT, XNOR_1_2_NAND2_NUM8_OUT, XNOR_1_3_NAND2_NUM8_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM8 (.ZN (XNOR_1_1_NAND2_NUM8_OUT), .A1 (N113), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM8 (.ZN (XNOR_1_2_NAND2_NUM8_OUT), .A1 (GND), .A2 (N120));
      NOR2_X1 XNOR_1_3_NAND2_NUM8 (.ZN (XNOR_1_3_NAND2_NUM8_OUT), .A1 (XNOR_1_1_NAND2_NUM8_OUT), .A2 (XNOR_1_2_NAND2_NUM8_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM8 (.ZN (N290), .A1 (XNOR_1_3_NAND2_NUM8_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM9_OUT, XNOR_1_2_NAND2_NUM9_OUT, XNOR_1_3_NAND2_NUM9_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM9 (.ZN (XNOR_1_1_NAND2_NUM9_OUT), .A1 (N127), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM9 (.ZN (XNOR_1_2_NAND2_NUM9_OUT), .A1 (GND), .A2 (N134));
      NOR2_X1 XNOR_1_3_NAND2_NUM9 (.ZN (XNOR_1_3_NAND2_NUM9_OUT), .A1 (XNOR_1_1_NAND2_NUM9_OUT), .A2 (XNOR_1_2_NAND2_NUM9_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM9 (.ZN (N293), .A1 (XNOR_1_3_NAND2_NUM9_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM10_OUT, XNOR_1_2_NAND2_NUM10_OUT, XNOR_1_3_NAND2_NUM10_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM10 (.ZN (XNOR_1_1_NAND2_NUM10_OUT), .A1 (N141), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM10 (.ZN (XNOR_1_2_NAND2_NUM10_OUT), .A1 (GND), .A2 (N148));
      NOR2_X1 XNOR_1_3_NAND2_NUM10 (.ZN (XNOR_1_3_NAND2_NUM10_OUT), .A1 (XNOR_1_1_NAND2_NUM10_OUT), .A2 (XNOR_1_2_NAND2_NUM10_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM10 (.ZN (N296), .A1 (XNOR_1_3_NAND2_NUM10_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM11_OUT, XNOR_1_2_NAND2_NUM11_OUT, XNOR_1_3_NAND2_NUM11_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM11 (.ZN (XNOR_1_1_NAND2_NUM11_OUT), .A1 (N155), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM11 (.ZN (XNOR_1_2_NAND2_NUM11_OUT), .A1 (GND), .A2 (N162));
      NOR2_X1 XNOR_1_3_NAND2_NUM11 (.ZN (XNOR_1_3_NAND2_NUM11_OUT), .A1 (XNOR_1_1_NAND2_NUM11_OUT), .A2 (XNOR_1_2_NAND2_NUM11_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM11 (.ZN (N299), .A1 (XNOR_1_3_NAND2_NUM11_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM12_OUT, XNOR_1_2_NAND2_NUM12_OUT, XNOR_1_3_NAND2_NUM12_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM12 (.ZN (XNOR_1_1_NAND2_NUM12_OUT), .A1 (N169), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM12 (.ZN (XNOR_1_2_NAND2_NUM12_OUT), .A1 (GND), .A2 (N176));
      NOR2_X1 XNOR_1_3_NAND2_NUM12 (.ZN (XNOR_1_3_NAND2_NUM12_OUT), .A1 (XNOR_1_1_NAND2_NUM12_OUT), .A2 (XNOR_1_2_NAND2_NUM12_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM12 (.ZN (N302), .A1 (XNOR_1_3_NAND2_NUM12_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM13_OUT, XNOR_1_2_NAND2_NUM13_OUT, XNOR_1_3_NAND2_NUM13_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM13 (.ZN (XNOR_1_1_NAND2_NUM13_OUT), .A1 (N183), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM13 (.ZN (XNOR_1_2_NAND2_NUM13_OUT), .A1 (GND), .A2 (N190));
      NOR2_X1 XNOR_1_3_NAND2_NUM13 (.ZN (XNOR_1_3_NAND2_NUM13_OUT), .A1 (XNOR_1_1_NAND2_NUM13_OUT), .A2 (XNOR_1_2_NAND2_NUM13_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM13 (.ZN (N305), .A1 (XNOR_1_3_NAND2_NUM13_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM14_OUT, XNOR_1_2_NAND2_NUM14_OUT, XNOR_1_3_NAND2_NUM14_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM14 (.ZN (XNOR_1_1_NAND2_NUM14_OUT), .A1 (N197), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM14 (.ZN (XNOR_1_2_NAND2_NUM14_OUT), .A1 (GND), .A2 (N204));
      NOR2_X1 XNOR_1_3_NAND2_NUM14 (.ZN (XNOR_1_3_NAND2_NUM14_OUT), .A1 (XNOR_1_1_NAND2_NUM14_OUT), .A2 (XNOR_1_2_NAND2_NUM14_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM14 (.ZN (N308), .A1 (XNOR_1_3_NAND2_NUM14_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM15_OUT, XNOR_1_2_NAND2_NUM15_OUT, XNOR_1_3_NAND2_NUM15_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM15 (.ZN (XNOR_1_1_NAND2_NUM15_OUT), .A1 (N211), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM15 (.ZN (XNOR_1_2_NAND2_NUM15_OUT), .A1 (GND), .A2 (N218));
      NOR2_X1 XNOR_1_3_NAND2_NUM15 (.ZN (XNOR_1_3_NAND2_NUM15_OUT), .A1 (XNOR_1_1_NAND2_NUM15_OUT), .A2 (XNOR_1_2_NAND2_NUM15_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM15 (.ZN (N311), .A1 (XNOR_1_3_NAND2_NUM15_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM16_OUT, XNOR_1_2_NAND2_NUM16_OUT, XNOR_1_3_NAND2_NUM16_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM16 (.ZN (XNOR_1_1_NAND2_NUM16_OUT), .A1 (N1), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM16 (.ZN (XNOR_1_2_NAND2_NUM16_OUT), .A1 (GND), .A2 (N29));
      NOR2_X1 XNOR_1_3_NAND2_NUM16 (.ZN (XNOR_1_3_NAND2_NUM16_OUT), .A1 (XNOR_1_1_NAND2_NUM16_OUT), .A2 (XNOR_1_2_NAND2_NUM16_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM16 (.ZN (N314), .A1 (XNOR_1_3_NAND2_NUM16_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM17_OUT, XNOR_1_2_NAND2_NUM17_OUT, XNOR_1_3_NAND2_NUM17_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM17 (.ZN (XNOR_1_1_NAND2_NUM17_OUT), .A1 (N57), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM17 (.ZN (XNOR_1_2_NAND2_NUM17_OUT), .A1 (GND), .A2 (N85));
      NOR2_X1 XNOR_1_3_NAND2_NUM17 (.ZN (XNOR_1_3_NAND2_NUM17_OUT), .A1 (XNOR_1_1_NAND2_NUM17_OUT), .A2 (XNOR_1_2_NAND2_NUM17_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM17 (.ZN (N317), .A1 (XNOR_1_3_NAND2_NUM17_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM18_OUT, XNOR_1_2_NAND2_NUM18_OUT, XNOR_1_3_NAND2_NUM18_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM18 (.ZN (XNOR_1_1_NAND2_NUM18_OUT), .A1 (N8), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM18 (.ZN (XNOR_1_2_NAND2_NUM18_OUT), .A1 (GND), .A2 (N36));
      NOR2_X1 XNOR_1_3_NAND2_NUM18 (.ZN (XNOR_1_3_NAND2_NUM18_OUT), .A1 (XNOR_1_1_NAND2_NUM18_OUT), .A2 (XNOR_1_2_NAND2_NUM18_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM18 (.ZN (N320), .A1 (XNOR_1_3_NAND2_NUM18_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM19_OUT, XNOR_1_2_NAND2_NUM19_OUT, XNOR_1_3_NAND2_NUM19_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM19 (.ZN (XNOR_1_1_NAND2_NUM19_OUT), .A1 (N64), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM19 (.ZN (XNOR_1_2_NAND2_NUM19_OUT), .A1 (GND), .A2 (N92));
      NOR2_X1 XNOR_1_3_NAND2_NUM19 (.ZN (XNOR_1_3_NAND2_NUM19_OUT), .A1 (XNOR_1_1_NAND2_NUM19_OUT), .A2 (XNOR_1_2_NAND2_NUM19_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM19 (.ZN (N323), .A1 (XNOR_1_3_NAND2_NUM19_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM20_OUT, XNOR_1_2_NAND2_NUM20_OUT, XNOR_1_3_NAND2_NUM20_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM20 (.ZN (XNOR_1_1_NAND2_NUM20_OUT), .A1 (N15), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM20 (.ZN (XNOR_1_2_NAND2_NUM20_OUT), .A1 (GND), .A2 (N43));
      NOR2_X1 XNOR_1_3_NAND2_NUM20 (.ZN (XNOR_1_3_NAND2_NUM20_OUT), .A1 (XNOR_1_1_NAND2_NUM20_OUT), .A2 (XNOR_1_2_NAND2_NUM20_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM20 (.ZN (N326), .A1 (XNOR_1_3_NAND2_NUM20_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM21_OUT, XNOR_1_2_NAND2_NUM21_OUT, XNOR_1_3_NAND2_NUM21_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM21 (.ZN (XNOR_1_1_NAND2_NUM21_OUT), .A1 (N71), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM21 (.ZN (XNOR_1_2_NAND2_NUM21_OUT), .A1 (GND), .A2 (N99));
      NOR2_X1 XNOR_1_3_NAND2_NUM21 (.ZN (XNOR_1_3_NAND2_NUM21_OUT), .A1 (XNOR_1_1_NAND2_NUM21_OUT), .A2 (XNOR_1_2_NAND2_NUM21_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM21 (.ZN (N329), .A1 (XNOR_1_3_NAND2_NUM21_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM22_OUT, XNOR_1_2_NAND2_NUM22_OUT, XNOR_1_3_NAND2_NUM22_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM22 (.ZN (XNOR_1_1_NAND2_NUM22_OUT), .A1 (N22), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM22 (.ZN (XNOR_1_2_NAND2_NUM22_OUT), .A1 (GND), .A2 (N50));
      NOR2_X1 XNOR_1_3_NAND2_NUM22 (.ZN (XNOR_1_3_NAND2_NUM22_OUT), .A1 (XNOR_1_1_NAND2_NUM22_OUT), .A2 (XNOR_1_2_NAND2_NUM22_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM22 (.ZN (N332), .A1 (XNOR_1_3_NAND2_NUM22_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM23_OUT, XNOR_1_2_NAND2_NUM23_OUT, XNOR_1_3_NAND2_NUM23_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM23 (.ZN (XNOR_1_1_NAND2_NUM23_OUT), .A1 (N78), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM23 (.ZN (XNOR_1_2_NAND2_NUM23_OUT), .A1 (GND), .A2 (N106));
      NOR2_X1 XNOR_1_3_NAND2_NUM23 (.ZN (XNOR_1_3_NAND2_NUM23_OUT), .A1 (XNOR_1_1_NAND2_NUM23_OUT), .A2 (XNOR_1_2_NAND2_NUM23_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM23 (.ZN (N335), .A1 (XNOR_1_3_NAND2_NUM23_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM24_OUT, XNOR_1_2_NAND2_NUM24_OUT, XNOR_1_3_NAND2_NUM24_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM24 (.ZN (XNOR_1_1_NAND2_NUM24_OUT), .A1 (N113), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM24 (.ZN (XNOR_1_2_NAND2_NUM24_OUT), .A1 (GND), .A2 (N141));
      NOR2_X1 XNOR_1_3_NAND2_NUM24 (.ZN (XNOR_1_3_NAND2_NUM24_OUT), .A1 (XNOR_1_1_NAND2_NUM24_OUT), .A2 (XNOR_1_2_NAND2_NUM24_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM24 (.ZN (N338), .A1 (XNOR_1_3_NAND2_NUM24_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM25_OUT, XNOR_1_2_NAND2_NUM25_OUT, XNOR_1_3_NAND2_NUM25_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM25 (.ZN (XNOR_1_1_NAND2_NUM25_OUT), .A1 (N169), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM25 (.ZN (XNOR_1_2_NAND2_NUM25_OUT), .A1 (GND), .A2 (N197));
      NOR2_X1 XNOR_1_3_NAND2_NUM25 (.ZN (XNOR_1_3_NAND2_NUM25_OUT), .A1 (XNOR_1_1_NAND2_NUM25_OUT), .A2 (XNOR_1_2_NAND2_NUM25_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM25 (.ZN (N341), .A1 (XNOR_1_3_NAND2_NUM25_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM26_OUT, XNOR_1_2_NAND2_NUM26_OUT, XNOR_1_3_NAND2_NUM26_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM26 (.ZN (XNOR_1_1_NAND2_NUM26_OUT), .A1 (N120), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM26 (.ZN (XNOR_1_2_NAND2_NUM26_OUT), .A1 (GND), .A2 (N148));
      NOR2_X1 XNOR_1_3_NAND2_NUM26 (.ZN (XNOR_1_3_NAND2_NUM26_OUT), .A1 (XNOR_1_1_NAND2_NUM26_OUT), .A2 (XNOR_1_2_NAND2_NUM26_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM26 (.ZN (N344), .A1 (XNOR_1_3_NAND2_NUM26_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM27_OUT, XNOR_1_2_NAND2_NUM27_OUT, XNOR_1_3_NAND2_NUM27_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM27 (.ZN (XNOR_1_1_NAND2_NUM27_OUT), .A1 (N176), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM27 (.ZN (XNOR_1_2_NAND2_NUM27_OUT), .A1 (GND), .A2 (N204));
      NOR2_X1 XNOR_1_3_NAND2_NUM27 (.ZN (XNOR_1_3_NAND2_NUM27_OUT), .A1 (XNOR_1_1_NAND2_NUM27_OUT), .A2 (XNOR_1_2_NAND2_NUM27_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM27 (.ZN (N347), .A1 (XNOR_1_3_NAND2_NUM27_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM28_OUT, XNOR_1_2_NAND2_NUM28_OUT, XNOR_1_3_NAND2_NUM28_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM28 (.ZN (XNOR_1_1_NAND2_NUM28_OUT), .A1 (N127), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM28 (.ZN (XNOR_1_2_NAND2_NUM28_OUT), .A1 (GND), .A2 (N155));
      NOR2_X1 XNOR_1_3_NAND2_NUM28 (.ZN (XNOR_1_3_NAND2_NUM28_OUT), .A1 (XNOR_1_1_NAND2_NUM28_OUT), .A2 (XNOR_1_2_NAND2_NUM28_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM28 (.ZN (N350), .A1 (XNOR_1_3_NAND2_NUM28_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM29_OUT, XNOR_1_2_NAND2_NUM29_OUT, XNOR_1_3_NAND2_NUM29_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM29 (.ZN (XNOR_1_1_NAND2_NUM29_OUT), .A1 (N183), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM29 (.ZN (XNOR_1_2_NAND2_NUM29_OUT), .A1 (GND), .A2 (N211));
      NOR2_X1 XNOR_1_3_NAND2_NUM29 (.ZN (XNOR_1_3_NAND2_NUM29_OUT), .A1 (XNOR_1_1_NAND2_NUM29_OUT), .A2 (XNOR_1_2_NAND2_NUM29_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM29 (.ZN (N353), .A1 (XNOR_1_3_NAND2_NUM29_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM30_OUT, XNOR_1_2_NAND2_NUM30_OUT, XNOR_1_3_NAND2_NUM30_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM30 (.ZN (XNOR_1_1_NAND2_NUM30_OUT), .A1 (N134), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM30 (.ZN (XNOR_1_2_NAND2_NUM30_OUT), .A1 (GND), .A2 (N162));
      NOR2_X1 XNOR_1_3_NAND2_NUM30 (.ZN (XNOR_1_3_NAND2_NUM30_OUT), .A1 (XNOR_1_1_NAND2_NUM30_OUT), .A2 (XNOR_1_2_NAND2_NUM30_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM30 (.ZN (N356), .A1 (XNOR_1_3_NAND2_NUM30_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM31_OUT, XNOR_1_2_NAND2_NUM31_OUT, XNOR_1_3_NAND2_NUM31_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM31 (.ZN (XNOR_1_1_NAND2_NUM31_OUT), .A1 (N190), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM31 (.ZN (XNOR_1_2_NAND2_NUM31_OUT), .A1 (GND), .A2 (N218));
      NOR2_X1 XNOR_1_3_NAND2_NUM31 (.ZN (XNOR_1_3_NAND2_NUM31_OUT), .A1 (XNOR_1_1_NAND2_NUM31_OUT), .A2 (XNOR_1_2_NAND2_NUM31_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM31 (.ZN (N359), .A1 (XNOR_1_3_NAND2_NUM31_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM32_OUT, XNOR_1_2_NAND2_NUM32_OUT, XNOR_1_3_NAND2_NUM32_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM32 (.ZN (XNOR_1_1_NAND2_NUM32_OUT), .A1 (N1), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM32 (.ZN (XNOR_1_2_NAND2_NUM32_OUT), .A1 (GND), .A2 (N266));
      NOR2_X1 XNOR_1_3_NAND2_NUM32 (.ZN (XNOR_1_3_NAND2_NUM32_OUT), .A1 (XNOR_1_1_NAND2_NUM32_OUT), .A2 (XNOR_1_2_NAND2_NUM32_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM32 (.ZN (N362), .A1 (XNOR_1_3_NAND2_NUM32_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM33_OUT, XNOR_1_2_NAND2_NUM33_OUT, XNOR_1_3_NAND2_NUM33_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM33 (.ZN (XNOR_1_1_NAND2_NUM33_OUT), .A1 (N8), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM33 (.ZN (XNOR_1_2_NAND2_NUM33_OUT), .A1 (GND), .A2 (N266));
      NOR2_X1 XNOR_1_3_NAND2_NUM33 (.ZN (XNOR_1_3_NAND2_NUM33_OUT), .A1 (XNOR_1_1_NAND2_NUM33_OUT), .A2 (XNOR_1_2_NAND2_NUM33_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM33 (.ZN (N363), .A1 (XNOR_1_3_NAND2_NUM33_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM34_OUT, XNOR_1_2_NAND2_NUM34_OUT, XNOR_1_3_NAND2_NUM34_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM34 (.ZN (XNOR_1_1_NAND2_NUM34_OUT), .A1 (N15), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM34 (.ZN (XNOR_1_2_NAND2_NUM34_OUT), .A1 (GND), .A2 (N269));
      NOR2_X1 XNOR_1_3_NAND2_NUM34 (.ZN (XNOR_1_3_NAND2_NUM34_OUT), .A1 (XNOR_1_1_NAND2_NUM34_OUT), .A2 (XNOR_1_2_NAND2_NUM34_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM34 (.ZN (N364), .A1 (XNOR_1_3_NAND2_NUM34_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM35_OUT, XNOR_1_2_NAND2_NUM35_OUT, XNOR_1_3_NAND2_NUM35_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM35 (.ZN (XNOR_1_1_NAND2_NUM35_OUT), .A1 (N22), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM35 (.ZN (XNOR_1_2_NAND2_NUM35_OUT), .A1 (GND), .A2 (N269));
      NOR2_X1 XNOR_1_3_NAND2_NUM35 (.ZN (XNOR_1_3_NAND2_NUM35_OUT), .A1 (XNOR_1_1_NAND2_NUM35_OUT), .A2 (XNOR_1_2_NAND2_NUM35_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM35 (.ZN (N365), .A1 (XNOR_1_3_NAND2_NUM35_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM36_OUT, XNOR_1_2_NAND2_NUM36_OUT, XNOR_1_3_NAND2_NUM36_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM36 (.ZN (XNOR_1_1_NAND2_NUM36_OUT), .A1 (N29), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM36 (.ZN (XNOR_1_2_NAND2_NUM36_OUT), .A1 (GND), .A2 (N272));
      NOR2_X1 XNOR_1_3_NAND2_NUM36 (.ZN (XNOR_1_3_NAND2_NUM36_OUT), .A1 (XNOR_1_1_NAND2_NUM36_OUT), .A2 (XNOR_1_2_NAND2_NUM36_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM36 (.ZN (N366), .A1 (XNOR_1_3_NAND2_NUM36_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM37_OUT, XNOR_1_2_NAND2_NUM37_OUT, XNOR_1_3_NAND2_NUM37_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM37 (.ZN (XNOR_1_1_NAND2_NUM37_OUT), .A1 (N36), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM37 (.ZN (XNOR_1_2_NAND2_NUM37_OUT), .A1 (GND), .A2 (N272));
      NOR2_X1 XNOR_1_3_NAND2_NUM37 (.ZN (XNOR_1_3_NAND2_NUM37_OUT), .A1 (XNOR_1_1_NAND2_NUM37_OUT), .A2 (XNOR_1_2_NAND2_NUM37_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM37 (.ZN (N367), .A1 (XNOR_1_3_NAND2_NUM37_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM38_OUT, XNOR_1_2_NAND2_NUM38_OUT, XNOR_1_3_NAND2_NUM38_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM38 (.ZN (XNOR_1_1_NAND2_NUM38_OUT), .A1 (N43), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM38 (.ZN (XNOR_1_2_NAND2_NUM38_OUT), .A1 (GND), .A2 (N275));
      NOR2_X1 XNOR_1_3_NAND2_NUM38 (.ZN (XNOR_1_3_NAND2_NUM38_OUT), .A1 (XNOR_1_1_NAND2_NUM38_OUT), .A2 (XNOR_1_2_NAND2_NUM38_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM38 (.ZN (N368), .A1 (XNOR_1_3_NAND2_NUM38_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM39_OUT, XNOR_1_2_NAND2_NUM39_OUT, XNOR_1_3_NAND2_NUM39_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM39 (.ZN (XNOR_1_1_NAND2_NUM39_OUT), .A1 (N50), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM39 (.ZN (XNOR_1_2_NAND2_NUM39_OUT), .A1 (GND), .A2 (N275));
      NOR2_X1 XNOR_1_3_NAND2_NUM39 (.ZN (XNOR_1_3_NAND2_NUM39_OUT), .A1 (XNOR_1_1_NAND2_NUM39_OUT), .A2 (XNOR_1_2_NAND2_NUM39_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM39 (.ZN (N369), .A1 (XNOR_1_3_NAND2_NUM39_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM40_OUT, XNOR_1_2_NAND2_NUM40_OUT, XNOR_1_3_NAND2_NUM40_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM40 (.ZN (XNOR_1_1_NAND2_NUM40_OUT), .A1 (N57), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM40 (.ZN (XNOR_1_2_NAND2_NUM40_OUT), .A1 (GND), .A2 (N278));
      NOR2_X1 XNOR_1_3_NAND2_NUM40 (.ZN (XNOR_1_3_NAND2_NUM40_OUT), .A1 (XNOR_1_1_NAND2_NUM40_OUT), .A2 (XNOR_1_2_NAND2_NUM40_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM40 (.ZN (N370), .A1 (XNOR_1_3_NAND2_NUM40_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM41_OUT, XNOR_1_2_NAND2_NUM41_OUT, XNOR_1_3_NAND2_NUM41_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM41 (.ZN (XNOR_1_1_NAND2_NUM41_OUT), .A1 (N64), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM41 (.ZN (XNOR_1_2_NAND2_NUM41_OUT), .A1 (GND), .A2 (N278));
      NOR2_X1 XNOR_1_3_NAND2_NUM41 (.ZN (XNOR_1_3_NAND2_NUM41_OUT), .A1 (XNOR_1_1_NAND2_NUM41_OUT), .A2 (XNOR_1_2_NAND2_NUM41_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM41 (.ZN (N371), .A1 (XNOR_1_3_NAND2_NUM41_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM42_OUT, XNOR_1_2_NAND2_NUM42_OUT, XNOR_1_3_NAND2_NUM42_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM42 (.ZN (XNOR_1_1_NAND2_NUM42_OUT), .A1 (N71), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM42 (.ZN (XNOR_1_2_NAND2_NUM42_OUT), .A1 (GND), .A2 (N281));
      NOR2_X1 XNOR_1_3_NAND2_NUM42 (.ZN (XNOR_1_3_NAND2_NUM42_OUT), .A1 (XNOR_1_1_NAND2_NUM42_OUT), .A2 (XNOR_1_2_NAND2_NUM42_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM42 (.ZN (N372), .A1 (XNOR_1_3_NAND2_NUM42_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM43_OUT, XNOR_1_2_NAND2_NUM43_OUT, XNOR_1_3_NAND2_NUM43_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM43 (.ZN (XNOR_1_1_NAND2_NUM43_OUT), .A1 (N78), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM43 (.ZN (XNOR_1_2_NAND2_NUM43_OUT), .A1 (GND), .A2 (N281));
      NOR2_X1 XNOR_1_3_NAND2_NUM43 (.ZN (XNOR_1_3_NAND2_NUM43_OUT), .A1 (XNOR_1_1_NAND2_NUM43_OUT), .A2 (XNOR_1_2_NAND2_NUM43_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM43 (.ZN (N373), .A1 (XNOR_1_3_NAND2_NUM43_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM44_OUT, XNOR_1_2_NAND2_NUM44_OUT, XNOR_1_3_NAND2_NUM44_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM44 (.ZN (XNOR_1_1_NAND2_NUM44_OUT), .A1 (N85), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM44 (.ZN (XNOR_1_2_NAND2_NUM44_OUT), .A1 (GND), .A2 (N284));
      NOR2_X1 XNOR_1_3_NAND2_NUM44 (.ZN (XNOR_1_3_NAND2_NUM44_OUT), .A1 (XNOR_1_1_NAND2_NUM44_OUT), .A2 (XNOR_1_2_NAND2_NUM44_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM44 (.ZN (N374), .A1 (XNOR_1_3_NAND2_NUM44_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM45_OUT, XNOR_1_2_NAND2_NUM45_OUT, XNOR_1_3_NAND2_NUM45_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM45 (.ZN (XNOR_1_1_NAND2_NUM45_OUT), .A1 (N92), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM45 (.ZN (XNOR_1_2_NAND2_NUM45_OUT), .A1 (GND), .A2 (N284));
      NOR2_X1 XNOR_1_3_NAND2_NUM45 (.ZN (XNOR_1_3_NAND2_NUM45_OUT), .A1 (XNOR_1_1_NAND2_NUM45_OUT), .A2 (XNOR_1_2_NAND2_NUM45_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM45 (.ZN (N375), .A1 (XNOR_1_3_NAND2_NUM45_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM46_OUT, XNOR_1_2_NAND2_NUM46_OUT, XNOR_1_3_NAND2_NUM46_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM46 (.ZN (XNOR_1_1_NAND2_NUM46_OUT), .A1 (N99), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM46 (.ZN (XNOR_1_2_NAND2_NUM46_OUT), .A1 (GND), .A2 (N287));
      NOR2_X1 XNOR_1_3_NAND2_NUM46 (.ZN (XNOR_1_3_NAND2_NUM46_OUT), .A1 (XNOR_1_1_NAND2_NUM46_OUT), .A2 (XNOR_1_2_NAND2_NUM46_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM46 (.ZN (N376), .A1 (XNOR_1_3_NAND2_NUM46_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM47_OUT, XNOR_1_2_NAND2_NUM47_OUT, XNOR_1_3_NAND2_NUM47_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM47 (.ZN (XNOR_1_1_NAND2_NUM47_OUT), .A1 (N106), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM47 (.ZN (XNOR_1_2_NAND2_NUM47_OUT), .A1 (GND), .A2 (N287));
      NOR2_X1 XNOR_1_3_NAND2_NUM47 (.ZN (XNOR_1_3_NAND2_NUM47_OUT), .A1 (XNOR_1_1_NAND2_NUM47_OUT), .A2 (XNOR_1_2_NAND2_NUM47_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM47 (.ZN (N377), .A1 (XNOR_1_3_NAND2_NUM47_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM48_OUT, XNOR_1_2_NAND2_NUM48_OUT, XNOR_1_3_NAND2_NUM48_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM48 (.ZN (XNOR_1_1_NAND2_NUM48_OUT), .A1 (N113), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM48 (.ZN (XNOR_1_2_NAND2_NUM48_OUT), .A1 (GND), .A2 (N290));
      NOR2_X1 XNOR_1_3_NAND2_NUM48 (.ZN (XNOR_1_3_NAND2_NUM48_OUT), .A1 (XNOR_1_1_NAND2_NUM48_OUT), .A2 (XNOR_1_2_NAND2_NUM48_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM48 (.ZN (N378), .A1 (XNOR_1_3_NAND2_NUM48_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM49_OUT, XNOR_1_2_NAND2_NUM49_OUT, XNOR_1_3_NAND2_NUM49_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM49 (.ZN (XNOR_1_1_NAND2_NUM49_OUT), .A1 (N120), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM49 (.ZN (XNOR_1_2_NAND2_NUM49_OUT), .A1 (GND), .A2 (N290));
      NOR2_X1 XNOR_1_3_NAND2_NUM49 (.ZN (XNOR_1_3_NAND2_NUM49_OUT), .A1 (XNOR_1_1_NAND2_NUM49_OUT), .A2 (XNOR_1_2_NAND2_NUM49_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM49 (.ZN (N379), .A1 (XNOR_1_3_NAND2_NUM49_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM50_OUT, XNOR_1_2_NAND2_NUM50_OUT, XNOR_1_3_NAND2_NUM50_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM50 (.ZN (XNOR_1_1_NAND2_NUM50_OUT), .A1 (N127), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM50 (.ZN (XNOR_1_2_NAND2_NUM50_OUT), .A1 (GND), .A2 (N293));
      NOR2_X1 XNOR_1_3_NAND2_NUM50 (.ZN (XNOR_1_3_NAND2_NUM50_OUT), .A1 (XNOR_1_1_NAND2_NUM50_OUT), .A2 (XNOR_1_2_NAND2_NUM50_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM50 (.ZN (N380), .A1 (XNOR_1_3_NAND2_NUM50_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM51_OUT, XNOR_1_2_NAND2_NUM51_OUT, XNOR_1_3_NAND2_NUM51_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM51 (.ZN (XNOR_1_1_NAND2_NUM51_OUT), .A1 (N134), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM51 (.ZN (XNOR_1_2_NAND2_NUM51_OUT), .A1 (GND), .A2 (N293));
      NOR2_X1 XNOR_1_3_NAND2_NUM51 (.ZN (XNOR_1_3_NAND2_NUM51_OUT), .A1 (XNOR_1_1_NAND2_NUM51_OUT), .A2 (XNOR_1_2_NAND2_NUM51_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM51 (.ZN (N381), .A1 (XNOR_1_3_NAND2_NUM51_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM52_OUT, XNOR_1_2_NAND2_NUM52_OUT, XNOR_1_3_NAND2_NUM52_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM52 (.ZN (XNOR_1_1_NAND2_NUM52_OUT), .A1 (N141), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM52 (.ZN (XNOR_1_2_NAND2_NUM52_OUT), .A1 (GND), .A2 (N296));
      NOR2_X1 XNOR_1_3_NAND2_NUM52 (.ZN (XNOR_1_3_NAND2_NUM52_OUT), .A1 (XNOR_1_1_NAND2_NUM52_OUT), .A2 (XNOR_1_2_NAND2_NUM52_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM52 (.ZN (N382), .A1 (XNOR_1_3_NAND2_NUM52_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM53_OUT, XNOR_1_2_NAND2_NUM53_OUT, XNOR_1_3_NAND2_NUM53_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM53 (.ZN (XNOR_1_1_NAND2_NUM53_OUT), .A1 (N148), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM53 (.ZN (XNOR_1_2_NAND2_NUM53_OUT), .A1 (GND), .A2 (N296));
      NOR2_X1 XNOR_1_3_NAND2_NUM53 (.ZN (XNOR_1_3_NAND2_NUM53_OUT), .A1 (XNOR_1_1_NAND2_NUM53_OUT), .A2 (XNOR_1_2_NAND2_NUM53_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM53 (.ZN (N383), .A1 (XNOR_1_3_NAND2_NUM53_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM54_OUT, XNOR_1_2_NAND2_NUM54_OUT, XNOR_1_3_NAND2_NUM54_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM54 (.ZN (XNOR_1_1_NAND2_NUM54_OUT), .A1 (N155), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM54 (.ZN (XNOR_1_2_NAND2_NUM54_OUT), .A1 (GND), .A2 (N299));
      NOR2_X1 XNOR_1_3_NAND2_NUM54 (.ZN (XNOR_1_3_NAND2_NUM54_OUT), .A1 (XNOR_1_1_NAND2_NUM54_OUT), .A2 (XNOR_1_2_NAND2_NUM54_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM54 (.ZN (N384), .A1 (XNOR_1_3_NAND2_NUM54_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM55_OUT, XNOR_1_2_NAND2_NUM55_OUT, XNOR_1_3_NAND2_NUM55_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM55 (.ZN (XNOR_1_1_NAND2_NUM55_OUT), .A1 (N162), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM55 (.ZN (XNOR_1_2_NAND2_NUM55_OUT), .A1 (GND), .A2 (N299));
      NOR2_X1 XNOR_1_3_NAND2_NUM55 (.ZN (XNOR_1_3_NAND2_NUM55_OUT), .A1 (XNOR_1_1_NAND2_NUM55_OUT), .A2 (XNOR_1_2_NAND2_NUM55_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM55 (.ZN (N385), .A1 (XNOR_1_3_NAND2_NUM55_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM56_OUT, XNOR_1_2_NAND2_NUM56_OUT, XNOR_1_3_NAND2_NUM56_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM56 (.ZN (XNOR_1_1_NAND2_NUM56_OUT), .A1 (N169), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM56 (.ZN (XNOR_1_2_NAND2_NUM56_OUT), .A1 (GND), .A2 (N302));
      NOR2_X1 XNOR_1_3_NAND2_NUM56 (.ZN (XNOR_1_3_NAND2_NUM56_OUT), .A1 (XNOR_1_1_NAND2_NUM56_OUT), .A2 (XNOR_1_2_NAND2_NUM56_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM56 (.ZN (N386), .A1 (XNOR_1_3_NAND2_NUM56_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM57_OUT, XNOR_1_2_NAND2_NUM57_OUT, XNOR_1_3_NAND2_NUM57_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM57 (.ZN (XNOR_1_1_NAND2_NUM57_OUT), .A1 (N176), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM57 (.ZN (XNOR_1_2_NAND2_NUM57_OUT), .A1 (GND), .A2 (N302));
      NOR2_X1 XNOR_1_3_NAND2_NUM57 (.ZN (XNOR_1_3_NAND2_NUM57_OUT), .A1 (XNOR_1_1_NAND2_NUM57_OUT), .A2 (XNOR_1_2_NAND2_NUM57_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM57 (.ZN (N387), .A1 (XNOR_1_3_NAND2_NUM57_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM58_OUT, XNOR_1_2_NAND2_NUM58_OUT, XNOR_1_3_NAND2_NUM58_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM58 (.ZN (XNOR_1_1_NAND2_NUM58_OUT), .A1 (N183), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM58 (.ZN (XNOR_1_2_NAND2_NUM58_OUT), .A1 (GND), .A2 (N305));
      NOR2_X1 XNOR_1_3_NAND2_NUM58 (.ZN (XNOR_1_3_NAND2_NUM58_OUT), .A1 (XNOR_1_1_NAND2_NUM58_OUT), .A2 (XNOR_1_2_NAND2_NUM58_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM58 (.ZN (N388), .A1 (XNOR_1_3_NAND2_NUM58_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM59_OUT, XNOR_1_2_NAND2_NUM59_OUT, XNOR_1_3_NAND2_NUM59_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM59 (.ZN (XNOR_1_1_NAND2_NUM59_OUT), .A1 (N190), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM59 (.ZN (XNOR_1_2_NAND2_NUM59_OUT), .A1 (GND), .A2 (N305));
      NOR2_X1 XNOR_1_3_NAND2_NUM59 (.ZN (XNOR_1_3_NAND2_NUM59_OUT), .A1 (XNOR_1_1_NAND2_NUM59_OUT), .A2 (XNOR_1_2_NAND2_NUM59_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM59 (.ZN (N389), .A1 (XNOR_1_3_NAND2_NUM59_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM60_OUT, XNOR_1_2_NAND2_NUM60_OUT, XNOR_1_3_NAND2_NUM60_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM60 (.ZN (XNOR_1_1_NAND2_NUM60_OUT), .A1 (N197), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM60 (.ZN (XNOR_1_2_NAND2_NUM60_OUT), .A1 (GND), .A2 (N308));
      NOR2_X1 XNOR_1_3_NAND2_NUM60 (.ZN (XNOR_1_3_NAND2_NUM60_OUT), .A1 (XNOR_1_1_NAND2_NUM60_OUT), .A2 (XNOR_1_2_NAND2_NUM60_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM60 (.ZN (N390), .A1 (XNOR_1_3_NAND2_NUM60_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM61_OUT, XNOR_1_2_NAND2_NUM61_OUT, XNOR_1_3_NAND2_NUM61_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM61 (.ZN (XNOR_1_1_NAND2_NUM61_OUT), .A1 (N204), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM61 (.ZN (XNOR_1_2_NAND2_NUM61_OUT), .A1 (GND), .A2 (N308));
      NOR2_X1 XNOR_1_3_NAND2_NUM61 (.ZN (XNOR_1_3_NAND2_NUM61_OUT), .A1 (XNOR_1_1_NAND2_NUM61_OUT), .A2 (XNOR_1_2_NAND2_NUM61_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM61 (.ZN (N391), .A1 (XNOR_1_3_NAND2_NUM61_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM62_OUT, XNOR_1_2_NAND2_NUM62_OUT, XNOR_1_3_NAND2_NUM62_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM62 (.ZN (XNOR_1_1_NAND2_NUM62_OUT), .A1 (N211), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM62 (.ZN (XNOR_1_2_NAND2_NUM62_OUT), .A1 (GND), .A2 (N311));
      NOR2_X1 XNOR_1_3_NAND2_NUM62 (.ZN (XNOR_1_3_NAND2_NUM62_OUT), .A1 (XNOR_1_1_NAND2_NUM62_OUT), .A2 (XNOR_1_2_NAND2_NUM62_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM62 (.ZN (N392), .A1 (XNOR_1_3_NAND2_NUM62_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM63_OUT, XNOR_1_2_NAND2_NUM63_OUT, XNOR_1_3_NAND2_NUM63_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM63 (.ZN (XNOR_1_1_NAND2_NUM63_OUT), .A1 (N218), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM63 (.ZN (XNOR_1_2_NAND2_NUM63_OUT), .A1 (GND), .A2 (N311));
      NOR2_X1 XNOR_1_3_NAND2_NUM63 (.ZN (XNOR_1_3_NAND2_NUM63_OUT), .A1 (XNOR_1_1_NAND2_NUM63_OUT), .A2 (XNOR_1_2_NAND2_NUM63_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM63 (.ZN (N393), .A1 (XNOR_1_3_NAND2_NUM63_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM64_OUT, XNOR_1_2_NAND2_NUM64_OUT, XNOR_1_3_NAND2_NUM64_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM64 (.ZN (XNOR_1_1_NAND2_NUM64_OUT), .A1 (N1), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM64 (.ZN (XNOR_1_2_NAND2_NUM64_OUT), .A1 (GND), .A2 (N314));
      NOR2_X1 XNOR_1_3_NAND2_NUM64 (.ZN (XNOR_1_3_NAND2_NUM64_OUT), .A1 (XNOR_1_1_NAND2_NUM64_OUT), .A2 (XNOR_1_2_NAND2_NUM64_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM64 (.ZN (N394), .A1 (XNOR_1_3_NAND2_NUM64_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM65_OUT, XNOR_1_2_NAND2_NUM65_OUT, XNOR_1_3_NAND2_NUM65_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM65 (.ZN (XNOR_1_1_NAND2_NUM65_OUT), .A1 (N29), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM65 (.ZN (XNOR_1_2_NAND2_NUM65_OUT), .A1 (GND), .A2 (N314));
      NOR2_X1 XNOR_1_3_NAND2_NUM65 (.ZN (XNOR_1_3_NAND2_NUM65_OUT), .A1 (XNOR_1_1_NAND2_NUM65_OUT), .A2 (XNOR_1_2_NAND2_NUM65_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM65 (.ZN (N395), .A1 (XNOR_1_3_NAND2_NUM65_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM66_OUT, XNOR_1_2_NAND2_NUM66_OUT, XNOR_1_3_NAND2_NUM66_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM66 (.ZN (XNOR_1_1_NAND2_NUM66_OUT), .A1 (N57), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM66 (.ZN (XNOR_1_2_NAND2_NUM66_OUT), .A1 (GND), .A2 (N317));
      NOR2_X1 XNOR_1_3_NAND2_NUM66 (.ZN (XNOR_1_3_NAND2_NUM66_OUT), .A1 (XNOR_1_1_NAND2_NUM66_OUT), .A2 (XNOR_1_2_NAND2_NUM66_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM66 (.ZN (N396), .A1 (XNOR_1_3_NAND2_NUM66_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM67_OUT, XNOR_1_2_NAND2_NUM67_OUT, XNOR_1_3_NAND2_NUM67_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM67 (.ZN (XNOR_1_1_NAND2_NUM67_OUT), .A1 (N85), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM67 (.ZN (XNOR_1_2_NAND2_NUM67_OUT), .A1 (GND), .A2 (N317));
      NOR2_X1 XNOR_1_3_NAND2_NUM67 (.ZN (XNOR_1_3_NAND2_NUM67_OUT), .A1 (XNOR_1_1_NAND2_NUM67_OUT), .A2 (XNOR_1_2_NAND2_NUM67_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM67 (.ZN (N397), .A1 (XNOR_1_3_NAND2_NUM67_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM68_OUT, XNOR_1_2_NAND2_NUM68_OUT, XNOR_1_3_NAND2_NUM68_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM68 (.ZN (XNOR_1_1_NAND2_NUM68_OUT), .A1 (N8), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM68 (.ZN (XNOR_1_2_NAND2_NUM68_OUT), .A1 (GND), .A2 (N320));
      NOR2_X1 XNOR_1_3_NAND2_NUM68 (.ZN (XNOR_1_3_NAND2_NUM68_OUT), .A1 (XNOR_1_1_NAND2_NUM68_OUT), .A2 (XNOR_1_2_NAND2_NUM68_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM68 (.ZN (N398), .A1 (XNOR_1_3_NAND2_NUM68_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM69_OUT, XNOR_1_2_NAND2_NUM69_OUT, XNOR_1_3_NAND2_NUM69_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM69 (.ZN (XNOR_1_1_NAND2_NUM69_OUT), .A1 (N36), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM69 (.ZN (XNOR_1_2_NAND2_NUM69_OUT), .A1 (GND), .A2 (N320));
      NOR2_X1 XNOR_1_3_NAND2_NUM69 (.ZN (XNOR_1_3_NAND2_NUM69_OUT), .A1 (XNOR_1_1_NAND2_NUM69_OUT), .A2 (XNOR_1_2_NAND2_NUM69_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM69 (.ZN (N399), .A1 (XNOR_1_3_NAND2_NUM69_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM70_OUT, XNOR_1_2_NAND2_NUM70_OUT, XNOR_1_3_NAND2_NUM70_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM70 (.ZN (XNOR_1_1_NAND2_NUM70_OUT), .A1 (N64), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM70 (.ZN (XNOR_1_2_NAND2_NUM70_OUT), .A1 (GND), .A2 (N323));
      NOR2_X1 XNOR_1_3_NAND2_NUM70 (.ZN (XNOR_1_3_NAND2_NUM70_OUT), .A1 (XNOR_1_1_NAND2_NUM70_OUT), .A2 (XNOR_1_2_NAND2_NUM70_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM70 (.ZN (N400), .A1 (XNOR_1_3_NAND2_NUM70_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM71_OUT, XNOR_1_2_NAND2_NUM71_OUT, XNOR_1_3_NAND2_NUM71_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM71 (.ZN (XNOR_1_1_NAND2_NUM71_OUT), .A1 (N92), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM71 (.ZN (XNOR_1_2_NAND2_NUM71_OUT), .A1 (GND), .A2 (N323));
      NOR2_X1 XNOR_1_3_NAND2_NUM71 (.ZN (XNOR_1_3_NAND2_NUM71_OUT), .A1 (XNOR_1_1_NAND2_NUM71_OUT), .A2 (XNOR_1_2_NAND2_NUM71_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM71 (.ZN (N401), .A1 (XNOR_1_3_NAND2_NUM71_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM72_OUT, XNOR_1_2_NAND2_NUM72_OUT, XNOR_1_3_NAND2_NUM72_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM72 (.ZN (XNOR_1_1_NAND2_NUM72_OUT), .A1 (N15), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM72 (.ZN (XNOR_1_2_NAND2_NUM72_OUT), .A1 (GND), .A2 (N326));
      NOR2_X1 XNOR_1_3_NAND2_NUM72 (.ZN (XNOR_1_3_NAND2_NUM72_OUT), .A1 (XNOR_1_1_NAND2_NUM72_OUT), .A2 (XNOR_1_2_NAND2_NUM72_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM72 (.ZN (N402), .A1 (XNOR_1_3_NAND2_NUM72_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM73_OUT, XNOR_1_2_NAND2_NUM73_OUT, XNOR_1_3_NAND2_NUM73_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM73 (.ZN (XNOR_1_1_NAND2_NUM73_OUT), .A1 (N43), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM73 (.ZN (XNOR_1_2_NAND2_NUM73_OUT), .A1 (GND), .A2 (N326));
      NOR2_X1 XNOR_1_3_NAND2_NUM73 (.ZN (XNOR_1_3_NAND2_NUM73_OUT), .A1 (XNOR_1_1_NAND2_NUM73_OUT), .A2 (XNOR_1_2_NAND2_NUM73_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM73 (.ZN (N403), .A1 (XNOR_1_3_NAND2_NUM73_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM74_OUT, XNOR_1_2_NAND2_NUM74_OUT, XNOR_1_3_NAND2_NUM74_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM74 (.ZN (XNOR_1_1_NAND2_NUM74_OUT), .A1 (N71), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM74 (.ZN (XNOR_1_2_NAND2_NUM74_OUT), .A1 (GND), .A2 (N329));
      NOR2_X1 XNOR_1_3_NAND2_NUM74 (.ZN (XNOR_1_3_NAND2_NUM74_OUT), .A1 (XNOR_1_1_NAND2_NUM74_OUT), .A2 (XNOR_1_2_NAND2_NUM74_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM74 (.ZN (N404), .A1 (XNOR_1_3_NAND2_NUM74_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM75_OUT, XNOR_1_2_NAND2_NUM75_OUT, XNOR_1_3_NAND2_NUM75_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM75 (.ZN (XNOR_1_1_NAND2_NUM75_OUT), .A1 (N99), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM75 (.ZN (XNOR_1_2_NAND2_NUM75_OUT), .A1 (GND), .A2 (N329));
      NOR2_X1 XNOR_1_3_NAND2_NUM75 (.ZN (XNOR_1_3_NAND2_NUM75_OUT), .A1 (XNOR_1_1_NAND2_NUM75_OUT), .A2 (XNOR_1_2_NAND2_NUM75_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM75 (.ZN (N405), .A1 (XNOR_1_3_NAND2_NUM75_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM76_OUT, XNOR_1_2_NAND2_NUM76_OUT, XNOR_1_3_NAND2_NUM76_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM76 (.ZN (XNOR_1_1_NAND2_NUM76_OUT), .A1 (N22), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM76 (.ZN (XNOR_1_2_NAND2_NUM76_OUT), .A1 (GND), .A2 (N332));
      NOR2_X1 XNOR_1_3_NAND2_NUM76 (.ZN (XNOR_1_3_NAND2_NUM76_OUT), .A1 (XNOR_1_1_NAND2_NUM76_OUT), .A2 (XNOR_1_2_NAND2_NUM76_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM76 (.ZN (N406), .A1 (XNOR_1_3_NAND2_NUM76_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM77_OUT, XNOR_1_2_NAND2_NUM77_OUT, XNOR_1_3_NAND2_NUM77_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM77 (.ZN (XNOR_1_1_NAND2_NUM77_OUT), .A1 (N50), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM77 (.ZN (XNOR_1_2_NAND2_NUM77_OUT), .A1 (GND), .A2 (N332));
      NOR2_X1 XNOR_1_3_NAND2_NUM77 (.ZN (XNOR_1_3_NAND2_NUM77_OUT), .A1 (XNOR_1_1_NAND2_NUM77_OUT), .A2 (XNOR_1_2_NAND2_NUM77_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM77 (.ZN (N407), .A1 (XNOR_1_3_NAND2_NUM77_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM78_OUT, XNOR_1_2_NAND2_NUM78_OUT, XNOR_1_3_NAND2_NUM78_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM78 (.ZN (XNOR_1_1_NAND2_NUM78_OUT), .A1 (N78), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM78 (.ZN (XNOR_1_2_NAND2_NUM78_OUT), .A1 (GND), .A2 (N335));
      NOR2_X1 XNOR_1_3_NAND2_NUM78 (.ZN (XNOR_1_3_NAND2_NUM78_OUT), .A1 (XNOR_1_1_NAND2_NUM78_OUT), .A2 (XNOR_1_2_NAND2_NUM78_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM78 (.ZN (N408), .A1 (XNOR_1_3_NAND2_NUM78_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM79_OUT, XNOR_1_2_NAND2_NUM79_OUT, XNOR_1_3_NAND2_NUM79_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM79 (.ZN (XNOR_1_1_NAND2_NUM79_OUT), .A1 (N106), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM79 (.ZN (XNOR_1_2_NAND2_NUM79_OUT), .A1 (GND), .A2 (N335));
      NOR2_X1 XNOR_1_3_NAND2_NUM79 (.ZN (XNOR_1_3_NAND2_NUM79_OUT), .A1 (XNOR_1_1_NAND2_NUM79_OUT), .A2 (XNOR_1_2_NAND2_NUM79_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM79 (.ZN (N409), .A1 (XNOR_1_3_NAND2_NUM79_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM80_OUT, XNOR_1_2_NAND2_NUM80_OUT, XNOR_1_3_NAND2_NUM80_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM80 (.ZN (XNOR_1_1_NAND2_NUM80_OUT), .A1 (N113), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM80 (.ZN (XNOR_1_2_NAND2_NUM80_OUT), .A1 (GND), .A2 (N338));
      NOR2_X1 XNOR_1_3_NAND2_NUM80 (.ZN (XNOR_1_3_NAND2_NUM80_OUT), .A1 (XNOR_1_1_NAND2_NUM80_OUT), .A2 (XNOR_1_2_NAND2_NUM80_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM80 (.ZN (N410), .A1 (XNOR_1_3_NAND2_NUM80_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM81_OUT, XNOR_1_2_NAND2_NUM81_OUT, XNOR_1_3_NAND2_NUM81_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM81 (.ZN (XNOR_1_1_NAND2_NUM81_OUT), .A1 (N141), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM81 (.ZN (XNOR_1_2_NAND2_NUM81_OUT), .A1 (GND), .A2 (N338));
      NOR2_X1 XNOR_1_3_NAND2_NUM81 (.ZN (XNOR_1_3_NAND2_NUM81_OUT), .A1 (XNOR_1_1_NAND2_NUM81_OUT), .A2 (XNOR_1_2_NAND2_NUM81_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM81 (.ZN (N411), .A1 (XNOR_1_3_NAND2_NUM81_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM82_OUT, XNOR_1_2_NAND2_NUM82_OUT, XNOR_1_3_NAND2_NUM82_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM82 (.ZN (XNOR_1_1_NAND2_NUM82_OUT), .A1 (N169), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM82 (.ZN (XNOR_1_2_NAND2_NUM82_OUT), .A1 (GND), .A2 (N341));
      NOR2_X1 XNOR_1_3_NAND2_NUM82 (.ZN (XNOR_1_3_NAND2_NUM82_OUT), .A1 (XNOR_1_1_NAND2_NUM82_OUT), .A2 (XNOR_1_2_NAND2_NUM82_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM82 (.ZN (N412), .A1 (XNOR_1_3_NAND2_NUM82_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM83_OUT, XNOR_1_2_NAND2_NUM83_OUT, XNOR_1_3_NAND2_NUM83_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM83 (.ZN (XNOR_1_1_NAND2_NUM83_OUT), .A1 (N197), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM83 (.ZN (XNOR_1_2_NAND2_NUM83_OUT), .A1 (GND), .A2 (N341));
      NOR2_X1 XNOR_1_3_NAND2_NUM83 (.ZN (XNOR_1_3_NAND2_NUM83_OUT), .A1 (XNOR_1_1_NAND2_NUM83_OUT), .A2 (XNOR_1_2_NAND2_NUM83_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM83 (.ZN (N413), .A1 (XNOR_1_3_NAND2_NUM83_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM84_OUT, XNOR_1_2_NAND2_NUM84_OUT, XNOR_1_3_NAND2_NUM84_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM84 (.ZN (XNOR_1_1_NAND2_NUM84_OUT), .A1 (N120), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM84 (.ZN (XNOR_1_2_NAND2_NUM84_OUT), .A1 (GND), .A2 (N344));
      NOR2_X1 XNOR_1_3_NAND2_NUM84 (.ZN (XNOR_1_3_NAND2_NUM84_OUT), .A1 (XNOR_1_1_NAND2_NUM84_OUT), .A2 (XNOR_1_2_NAND2_NUM84_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM84 (.ZN (N414), .A1 (XNOR_1_3_NAND2_NUM84_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM85_OUT, XNOR_1_2_NAND2_NUM85_OUT, XNOR_1_3_NAND2_NUM85_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM85 (.ZN (XNOR_1_1_NAND2_NUM85_OUT), .A1 (N148), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM85 (.ZN (XNOR_1_2_NAND2_NUM85_OUT), .A1 (GND), .A2 (N344));
      NOR2_X1 XNOR_1_3_NAND2_NUM85 (.ZN (XNOR_1_3_NAND2_NUM85_OUT), .A1 (XNOR_1_1_NAND2_NUM85_OUT), .A2 (XNOR_1_2_NAND2_NUM85_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM85 (.ZN (N415), .A1 (XNOR_1_3_NAND2_NUM85_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM86_OUT, XNOR_1_2_NAND2_NUM86_OUT, XNOR_1_3_NAND2_NUM86_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM86 (.ZN (XNOR_1_1_NAND2_NUM86_OUT), .A1 (N176), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM86 (.ZN (XNOR_1_2_NAND2_NUM86_OUT), .A1 (GND), .A2 (N347));
      NOR2_X1 XNOR_1_3_NAND2_NUM86 (.ZN (XNOR_1_3_NAND2_NUM86_OUT), .A1 (XNOR_1_1_NAND2_NUM86_OUT), .A2 (XNOR_1_2_NAND2_NUM86_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM86 (.ZN (N416), .A1 (XNOR_1_3_NAND2_NUM86_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM87_OUT, XNOR_1_2_NAND2_NUM87_OUT, XNOR_1_3_NAND2_NUM87_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM87 (.ZN (XNOR_1_1_NAND2_NUM87_OUT), .A1 (N204), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM87 (.ZN (XNOR_1_2_NAND2_NUM87_OUT), .A1 (GND), .A2 (N347));
      NOR2_X1 XNOR_1_3_NAND2_NUM87 (.ZN (XNOR_1_3_NAND2_NUM87_OUT), .A1 (XNOR_1_1_NAND2_NUM87_OUT), .A2 (XNOR_1_2_NAND2_NUM87_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM87 (.ZN (N417), .A1 (XNOR_1_3_NAND2_NUM87_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM88_OUT, XNOR_1_2_NAND2_NUM88_OUT, XNOR_1_3_NAND2_NUM88_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM88 (.ZN (XNOR_1_1_NAND2_NUM88_OUT), .A1 (N127), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM88 (.ZN (XNOR_1_2_NAND2_NUM88_OUT), .A1 (GND), .A2 (N350));
      NOR2_X1 XNOR_1_3_NAND2_NUM88 (.ZN (XNOR_1_3_NAND2_NUM88_OUT), .A1 (XNOR_1_1_NAND2_NUM88_OUT), .A2 (XNOR_1_2_NAND2_NUM88_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM88 (.ZN (N418), .A1 (XNOR_1_3_NAND2_NUM88_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM89_OUT, XNOR_1_2_NAND2_NUM89_OUT, XNOR_1_3_NAND2_NUM89_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM89 (.ZN (XNOR_1_1_NAND2_NUM89_OUT), .A1 (N155), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM89 (.ZN (XNOR_1_2_NAND2_NUM89_OUT), .A1 (GND), .A2 (N350));
      NOR2_X1 XNOR_1_3_NAND2_NUM89 (.ZN (XNOR_1_3_NAND2_NUM89_OUT), .A1 (XNOR_1_1_NAND2_NUM89_OUT), .A2 (XNOR_1_2_NAND2_NUM89_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM89 (.ZN (N419), .A1 (XNOR_1_3_NAND2_NUM89_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM90_OUT, XNOR_1_2_NAND2_NUM90_OUT, XNOR_1_3_NAND2_NUM90_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM90 (.ZN (XNOR_1_1_NAND2_NUM90_OUT), .A1 (N183), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM90 (.ZN (XNOR_1_2_NAND2_NUM90_OUT), .A1 (GND), .A2 (N353));
      NOR2_X1 XNOR_1_3_NAND2_NUM90 (.ZN (XNOR_1_3_NAND2_NUM90_OUT), .A1 (XNOR_1_1_NAND2_NUM90_OUT), .A2 (XNOR_1_2_NAND2_NUM90_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM90 (.ZN (N420), .A1 (XNOR_1_3_NAND2_NUM90_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM91_OUT, XNOR_1_2_NAND2_NUM91_OUT, XNOR_1_3_NAND2_NUM91_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM91 (.ZN (XNOR_1_1_NAND2_NUM91_OUT), .A1 (N211), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM91 (.ZN (XNOR_1_2_NAND2_NUM91_OUT), .A1 (GND), .A2 (N353));
      NOR2_X1 XNOR_1_3_NAND2_NUM91 (.ZN (XNOR_1_3_NAND2_NUM91_OUT), .A1 (XNOR_1_1_NAND2_NUM91_OUT), .A2 (XNOR_1_2_NAND2_NUM91_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM91 (.ZN (N421), .A1 (XNOR_1_3_NAND2_NUM91_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM92_OUT, XNOR_1_2_NAND2_NUM92_OUT, XNOR_1_3_NAND2_NUM92_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM92 (.ZN (XNOR_1_1_NAND2_NUM92_OUT), .A1 (N134), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM92 (.ZN (XNOR_1_2_NAND2_NUM92_OUT), .A1 (GND), .A2 (N356));
      NOR2_X1 XNOR_1_3_NAND2_NUM92 (.ZN (XNOR_1_3_NAND2_NUM92_OUT), .A1 (XNOR_1_1_NAND2_NUM92_OUT), .A2 (XNOR_1_2_NAND2_NUM92_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM92 (.ZN (N422), .A1 (XNOR_1_3_NAND2_NUM92_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM93_OUT, XNOR_1_2_NAND2_NUM93_OUT, XNOR_1_3_NAND2_NUM93_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM93 (.ZN (XNOR_1_1_NAND2_NUM93_OUT), .A1 (N162), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM93 (.ZN (XNOR_1_2_NAND2_NUM93_OUT), .A1 (GND), .A2 (N356));
      NOR2_X1 XNOR_1_3_NAND2_NUM93 (.ZN (XNOR_1_3_NAND2_NUM93_OUT), .A1 (XNOR_1_1_NAND2_NUM93_OUT), .A2 (XNOR_1_2_NAND2_NUM93_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM93 (.ZN (N423), .A1 (XNOR_1_3_NAND2_NUM93_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM94_OUT, XNOR_1_2_NAND2_NUM94_OUT, XNOR_1_3_NAND2_NUM94_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM94 (.ZN (XNOR_1_1_NAND2_NUM94_OUT), .A1 (N190), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM94 (.ZN (XNOR_1_2_NAND2_NUM94_OUT), .A1 (GND), .A2 (N359));
      NOR2_X1 XNOR_1_3_NAND2_NUM94 (.ZN (XNOR_1_3_NAND2_NUM94_OUT), .A1 (XNOR_1_1_NAND2_NUM94_OUT), .A2 (XNOR_1_2_NAND2_NUM94_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM94 (.ZN (N424), .A1 (XNOR_1_3_NAND2_NUM94_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM95_OUT, XNOR_1_2_NAND2_NUM95_OUT, XNOR_1_3_NAND2_NUM95_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM95 (.ZN (XNOR_1_1_NAND2_NUM95_OUT), .A1 (N218), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM95 (.ZN (XNOR_1_2_NAND2_NUM95_OUT), .A1 (GND), .A2 (N359));
      NOR2_X1 XNOR_1_3_NAND2_NUM95 (.ZN (XNOR_1_3_NAND2_NUM95_OUT), .A1 (XNOR_1_1_NAND2_NUM95_OUT), .A2 (XNOR_1_2_NAND2_NUM95_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM95 (.ZN (N425), .A1 (XNOR_1_3_NAND2_NUM95_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM96_OUT, XNOR_1_2_NAND2_NUM96_OUT, XNOR_1_3_NAND2_NUM96_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM96 (.ZN (XNOR_1_1_NAND2_NUM96_OUT), .A1 (N362), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM96 (.ZN (XNOR_1_2_NAND2_NUM96_OUT), .A1 (GND), .A2 (N363));
      NOR2_X1 XNOR_1_3_NAND2_NUM96 (.ZN (XNOR_1_3_NAND2_NUM96_OUT), .A1 (XNOR_1_1_NAND2_NUM96_OUT), .A2 (XNOR_1_2_NAND2_NUM96_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM96 (.ZN (N426), .A1 (XNOR_1_3_NAND2_NUM96_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM97_OUT, XNOR_1_2_NAND2_NUM97_OUT, XNOR_1_3_NAND2_NUM97_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM97 (.ZN (XNOR_1_1_NAND2_NUM97_OUT), .A1 (N364), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM97 (.ZN (XNOR_1_2_NAND2_NUM97_OUT), .A1 (GND), .A2 (N365));
      NOR2_X1 XNOR_1_3_NAND2_NUM97 (.ZN (XNOR_1_3_NAND2_NUM97_OUT), .A1 (XNOR_1_1_NAND2_NUM97_OUT), .A2 (XNOR_1_2_NAND2_NUM97_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM97 (.ZN (N429), .A1 (XNOR_1_3_NAND2_NUM97_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM98_OUT, XNOR_1_2_NAND2_NUM98_OUT, XNOR_1_3_NAND2_NUM98_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM98 (.ZN (XNOR_1_1_NAND2_NUM98_OUT), .A1 (N366), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM98 (.ZN (XNOR_1_2_NAND2_NUM98_OUT), .A1 (GND), .A2 (N367));
      NOR2_X1 XNOR_1_3_NAND2_NUM98 (.ZN (XNOR_1_3_NAND2_NUM98_OUT), .A1 (XNOR_1_1_NAND2_NUM98_OUT), .A2 (XNOR_1_2_NAND2_NUM98_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM98 (.ZN (N432), .A1 (XNOR_1_3_NAND2_NUM98_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM99_OUT, XNOR_1_2_NAND2_NUM99_OUT, XNOR_1_3_NAND2_NUM99_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM99 (.ZN (XNOR_1_1_NAND2_NUM99_OUT), .A1 (N368), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM99 (.ZN (XNOR_1_2_NAND2_NUM99_OUT), .A1 (GND), .A2 (N369));
      NOR2_X1 XNOR_1_3_NAND2_NUM99 (.ZN (XNOR_1_3_NAND2_NUM99_OUT), .A1 (XNOR_1_1_NAND2_NUM99_OUT), .A2 (XNOR_1_2_NAND2_NUM99_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM99 (.ZN (N435), .A1 (XNOR_1_3_NAND2_NUM99_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM100_OUT, XNOR_1_2_NAND2_NUM100_OUT, XNOR_1_3_NAND2_NUM100_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM100 (.ZN (XNOR_1_1_NAND2_NUM100_OUT), .A1 (N370), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM100 (.ZN (XNOR_1_2_NAND2_NUM100_OUT), .A1 (GND), .A2 (N371));
      NOR2_X1 XNOR_1_3_NAND2_NUM100 (.ZN (XNOR_1_3_NAND2_NUM100_OUT), .A1 (XNOR_1_1_NAND2_NUM100_OUT), .A2 (XNOR_1_2_NAND2_NUM100_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM100 (.ZN (N438), .A1 (XNOR_1_3_NAND2_NUM100_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM101_OUT, XNOR_1_2_NAND2_NUM101_OUT, XNOR_1_3_NAND2_NUM101_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM101 (.ZN (XNOR_1_1_NAND2_NUM101_OUT), .A1 (N372), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM101 (.ZN (XNOR_1_2_NAND2_NUM101_OUT), .A1 (GND), .A2 (N373));
      NOR2_X1 XNOR_1_3_NAND2_NUM101 (.ZN (XNOR_1_3_NAND2_NUM101_OUT), .A1 (XNOR_1_1_NAND2_NUM101_OUT), .A2 (XNOR_1_2_NAND2_NUM101_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM101 (.ZN (N441), .A1 (XNOR_1_3_NAND2_NUM101_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM102_OUT, XNOR_1_2_NAND2_NUM102_OUT, XNOR_1_3_NAND2_NUM102_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM102 (.ZN (XNOR_1_1_NAND2_NUM102_OUT), .A1 (N374), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM102 (.ZN (XNOR_1_2_NAND2_NUM102_OUT), .A1 (GND), .A2 (N375));
      NOR2_X1 XNOR_1_3_NAND2_NUM102 (.ZN (XNOR_1_3_NAND2_NUM102_OUT), .A1 (XNOR_1_1_NAND2_NUM102_OUT), .A2 (XNOR_1_2_NAND2_NUM102_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM102 (.ZN (N444), .A1 (XNOR_1_3_NAND2_NUM102_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM103_OUT, XNOR_1_2_NAND2_NUM103_OUT, XNOR_1_3_NAND2_NUM103_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM103 (.ZN (XNOR_1_1_NAND2_NUM103_OUT), .A1 (N376), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM103 (.ZN (XNOR_1_2_NAND2_NUM103_OUT), .A1 (GND), .A2 (N377));
      NOR2_X1 XNOR_1_3_NAND2_NUM103 (.ZN (XNOR_1_3_NAND2_NUM103_OUT), .A1 (XNOR_1_1_NAND2_NUM103_OUT), .A2 (XNOR_1_2_NAND2_NUM103_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM103 (.ZN (N447), .A1 (XNOR_1_3_NAND2_NUM103_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM104_OUT, XNOR_1_2_NAND2_NUM104_OUT, XNOR_1_3_NAND2_NUM104_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM104 (.ZN (XNOR_1_1_NAND2_NUM104_OUT), .A1 (N378), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM104 (.ZN (XNOR_1_2_NAND2_NUM104_OUT), .A1 (GND), .A2 (N379));
      NOR2_X1 XNOR_1_3_NAND2_NUM104 (.ZN (XNOR_1_3_NAND2_NUM104_OUT), .A1 (XNOR_1_1_NAND2_NUM104_OUT), .A2 (XNOR_1_2_NAND2_NUM104_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM104 (.ZN (N450), .A1 (XNOR_1_3_NAND2_NUM104_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM105_OUT, XNOR_1_2_NAND2_NUM105_OUT, XNOR_1_3_NAND2_NUM105_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM105 (.ZN (XNOR_1_1_NAND2_NUM105_OUT), .A1 (N380), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM105 (.ZN (XNOR_1_2_NAND2_NUM105_OUT), .A1 (GND), .A2 (N381));
      NOR2_X1 XNOR_1_3_NAND2_NUM105 (.ZN (XNOR_1_3_NAND2_NUM105_OUT), .A1 (XNOR_1_1_NAND2_NUM105_OUT), .A2 (XNOR_1_2_NAND2_NUM105_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM105 (.ZN (N453), .A1 (XNOR_1_3_NAND2_NUM105_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM106_OUT, XNOR_1_2_NAND2_NUM106_OUT, XNOR_1_3_NAND2_NUM106_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM106 (.ZN (XNOR_1_1_NAND2_NUM106_OUT), .A1 (N382), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM106 (.ZN (XNOR_1_2_NAND2_NUM106_OUT), .A1 (GND), .A2 (N383));
      NOR2_X1 XNOR_1_3_NAND2_NUM106 (.ZN (XNOR_1_3_NAND2_NUM106_OUT), .A1 (XNOR_1_1_NAND2_NUM106_OUT), .A2 (XNOR_1_2_NAND2_NUM106_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM106 (.ZN (N456), .A1 (XNOR_1_3_NAND2_NUM106_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM107_OUT, XNOR_1_2_NAND2_NUM107_OUT, XNOR_1_3_NAND2_NUM107_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM107 (.ZN (XNOR_1_1_NAND2_NUM107_OUT), .A1 (N384), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM107 (.ZN (XNOR_1_2_NAND2_NUM107_OUT), .A1 (GND), .A2 (N385));
      NOR2_X1 XNOR_1_3_NAND2_NUM107 (.ZN (XNOR_1_3_NAND2_NUM107_OUT), .A1 (XNOR_1_1_NAND2_NUM107_OUT), .A2 (XNOR_1_2_NAND2_NUM107_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM107 (.ZN (N459), .A1 (XNOR_1_3_NAND2_NUM107_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM108_OUT, XNOR_1_2_NAND2_NUM108_OUT, XNOR_1_3_NAND2_NUM108_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM108 (.ZN (XNOR_1_1_NAND2_NUM108_OUT), .A1 (N386), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM108 (.ZN (XNOR_1_2_NAND2_NUM108_OUT), .A1 (GND), .A2 (N387));
      NOR2_X1 XNOR_1_3_NAND2_NUM108 (.ZN (XNOR_1_3_NAND2_NUM108_OUT), .A1 (XNOR_1_1_NAND2_NUM108_OUT), .A2 (XNOR_1_2_NAND2_NUM108_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM108 (.ZN (N462), .A1 (XNOR_1_3_NAND2_NUM108_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM109_OUT, XNOR_1_2_NAND2_NUM109_OUT, XNOR_1_3_NAND2_NUM109_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM109 (.ZN (XNOR_1_1_NAND2_NUM109_OUT), .A1 (N388), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM109 (.ZN (XNOR_1_2_NAND2_NUM109_OUT), .A1 (GND), .A2 (N389));
      NOR2_X1 XNOR_1_3_NAND2_NUM109 (.ZN (XNOR_1_3_NAND2_NUM109_OUT), .A1 (XNOR_1_1_NAND2_NUM109_OUT), .A2 (XNOR_1_2_NAND2_NUM109_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM109 (.ZN (N465), .A1 (XNOR_1_3_NAND2_NUM109_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM110_OUT, XNOR_1_2_NAND2_NUM110_OUT, XNOR_1_3_NAND2_NUM110_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM110 (.ZN (XNOR_1_1_NAND2_NUM110_OUT), .A1 (N390), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM110 (.ZN (XNOR_1_2_NAND2_NUM110_OUT), .A1 (GND), .A2 (N391));
      NOR2_X1 XNOR_1_3_NAND2_NUM110 (.ZN (XNOR_1_3_NAND2_NUM110_OUT), .A1 (XNOR_1_1_NAND2_NUM110_OUT), .A2 (XNOR_1_2_NAND2_NUM110_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM110 (.ZN (N468), .A1 (XNOR_1_3_NAND2_NUM110_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM111_OUT, XNOR_1_2_NAND2_NUM111_OUT, XNOR_1_3_NAND2_NUM111_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM111 (.ZN (XNOR_1_1_NAND2_NUM111_OUT), .A1 (N392), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM111 (.ZN (XNOR_1_2_NAND2_NUM111_OUT), .A1 (GND), .A2 (N393));
      NOR2_X1 XNOR_1_3_NAND2_NUM111 (.ZN (XNOR_1_3_NAND2_NUM111_OUT), .A1 (XNOR_1_1_NAND2_NUM111_OUT), .A2 (XNOR_1_2_NAND2_NUM111_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM111 (.ZN (N471), .A1 (XNOR_1_3_NAND2_NUM111_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM112_OUT, XNOR_1_2_NAND2_NUM112_OUT, XNOR_1_3_NAND2_NUM112_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM112 (.ZN (XNOR_1_1_NAND2_NUM112_OUT), .A1 (N394), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM112 (.ZN (XNOR_1_2_NAND2_NUM112_OUT), .A1 (GND), .A2 (N395));
      NOR2_X1 XNOR_1_3_NAND2_NUM112 (.ZN (XNOR_1_3_NAND2_NUM112_OUT), .A1 (XNOR_1_1_NAND2_NUM112_OUT), .A2 (XNOR_1_2_NAND2_NUM112_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM112 (.ZN (N474), .A1 (XNOR_1_3_NAND2_NUM112_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM113_OUT, XNOR_1_2_NAND2_NUM113_OUT, XNOR_1_3_NAND2_NUM113_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM113 (.ZN (XNOR_1_1_NAND2_NUM113_OUT), .A1 (N396), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM113 (.ZN (XNOR_1_2_NAND2_NUM113_OUT), .A1 (GND), .A2 (N397));
      NOR2_X1 XNOR_1_3_NAND2_NUM113 (.ZN (XNOR_1_3_NAND2_NUM113_OUT), .A1 (XNOR_1_1_NAND2_NUM113_OUT), .A2 (XNOR_1_2_NAND2_NUM113_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM113 (.ZN (N477), .A1 (XNOR_1_3_NAND2_NUM113_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM114_OUT, XNOR_1_2_NAND2_NUM114_OUT, XNOR_1_3_NAND2_NUM114_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM114 (.ZN (XNOR_1_1_NAND2_NUM114_OUT), .A1 (N398), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM114 (.ZN (XNOR_1_2_NAND2_NUM114_OUT), .A1 (GND), .A2 (N399));
      NOR2_X1 XNOR_1_3_NAND2_NUM114 (.ZN (XNOR_1_3_NAND2_NUM114_OUT), .A1 (XNOR_1_1_NAND2_NUM114_OUT), .A2 (XNOR_1_2_NAND2_NUM114_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM114 (.ZN (N480), .A1 (XNOR_1_3_NAND2_NUM114_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM115_OUT, XNOR_1_2_NAND2_NUM115_OUT, XNOR_1_3_NAND2_NUM115_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM115 (.ZN (XNOR_1_1_NAND2_NUM115_OUT), .A1 (N400), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM115 (.ZN (XNOR_1_2_NAND2_NUM115_OUT), .A1 (GND), .A2 (N401));
      NOR2_X1 XNOR_1_3_NAND2_NUM115 (.ZN (XNOR_1_3_NAND2_NUM115_OUT), .A1 (XNOR_1_1_NAND2_NUM115_OUT), .A2 (XNOR_1_2_NAND2_NUM115_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM115 (.ZN (N483), .A1 (XNOR_1_3_NAND2_NUM115_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM116_OUT, XNOR_1_2_NAND2_NUM116_OUT, XNOR_1_3_NAND2_NUM116_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM116 (.ZN (XNOR_1_1_NAND2_NUM116_OUT), .A1 (N402), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM116 (.ZN (XNOR_1_2_NAND2_NUM116_OUT), .A1 (GND), .A2 (N403));
      NOR2_X1 XNOR_1_3_NAND2_NUM116 (.ZN (XNOR_1_3_NAND2_NUM116_OUT), .A1 (XNOR_1_1_NAND2_NUM116_OUT), .A2 (XNOR_1_2_NAND2_NUM116_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM116 (.ZN (N486), .A1 (XNOR_1_3_NAND2_NUM116_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM117_OUT, XNOR_1_2_NAND2_NUM117_OUT, XNOR_1_3_NAND2_NUM117_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM117 (.ZN (XNOR_1_1_NAND2_NUM117_OUT), .A1 (N404), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM117 (.ZN (XNOR_1_2_NAND2_NUM117_OUT), .A1 (GND), .A2 (N405));
      NOR2_X1 XNOR_1_3_NAND2_NUM117 (.ZN (XNOR_1_3_NAND2_NUM117_OUT), .A1 (XNOR_1_1_NAND2_NUM117_OUT), .A2 (XNOR_1_2_NAND2_NUM117_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM117 (.ZN (N489), .A1 (XNOR_1_3_NAND2_NUM117_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM118_OUT, XNOR_1_2_NAND2_NUM118_OUT, XNOR_1_3_NAND2_NUM118_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM118 (.ZN (XNOR_1_1_NAND2_NUM118_OUT), .A1 (N406), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM118 (.ZN (XNOR_1_2_NAND2_NUM118_OUT), .A1 (GND), .A2 (N407));
      NOR2_X1 XNOR_1_3_NAND2_NUM118 (.ZN (XNOR_1_3_NAND2_NUM118_OUT), .A1 (XNOR_1_1_NAND2_NUM118_OUT), .A2 (XNOR_1_2_NAND2_NUM118_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM118 (.ZN (N492), .A1 (XNOR_1_3_NAND2_NUM118_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM119_OUT, XNOR_1_2_NAND2_NUM119_OUT, XNOR_1_3_NAND2_NUM119_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM119 (.ZN (XNOR_1_1_NAND2_NUM119_OUT), .A1 (N408), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM119 (.ZN (XNOR_1_2_NAND2_NUM119_OUT), .A1 (GND), .A2 (N409));
      NOR2_X1 XNOR_1_3_NAND2_NUM119 (.ZN (XNOR_1_3_NAND2_NUM119_OUT), .A1 (XNOR_1_1_NAND2_NUM119_OUT), .A2 (XNOR_1_2_NAND2_NUM119_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM119 (.ZN (N495), .A1 (XNOR_1_3_NAND2_NUM119_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM120_OUT, XNOR_1_2_NAND2_NUM120_OUT, XNOR_1_3_NAND2_NUM120_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM120 (.ZN (XNOR_1_1_NAND2_NUM120_OUT), .A1 (N410), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM120 (.ZN (XNOR_1_2_NAND2_NUM120_OUT), .A1 (GND), .A2 (N411));
      NOR2_X1 XNOR_1_3_NAND2_NUM120 (.ZN (XNOR_1_3_NAND2_NUM120_OUT), .A1 (XNOR_1_1_NAND2_NUM120_OUT), .A2 (XNOR_1_2_NAND2_NUM120_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM120 (.ZN (N498), .A1 (XNOR_1_3_NAND2_NUM120_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM121_OUT, XNOR_1_2_NAND2_NUM121_OUT, XNOR_1_3_NAND2_NUM121_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM121 (.ZN (XNOR_1_1_NAND2_NUM121_OUT), .A1 (N412), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM121 (.ZN (XNOR_1_2_NAND2_NUM121_OUT), .A1 (GND), .A2 (N413));
      NOR2_X1 XNOR_1_3_NAND2_NUM121 (.ZN (XNOR_1_3_NAND2_NUM121_OUT), .A1 (XNOR_1_1_NAND2_NUM121_OUT), .A2 (XNOR_1_2_NAND2_NUM121_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM121 (.ZN (N501), .A1 (XNOR_1_3_NAND2_NUM121_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM122_OUT, XNOR_1_2_NAND2_NUM122_OUT, XNOR_1_3_NAND2_NUM122_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM122 (.ZN (XNOR_1_1_NAND2_NUM122_OUT), .A1 (N414), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM122 (.ZN (XNOR_1_2_NAND2_NUM122_OUT), .A1 (GND), .A2 (N415));
      NOR2_X1 XNOR_1_3_NAND2_NUM122 (.ZN (XNOR_1_3_NAND2_NUM122_OUT), .A1 (XNOR_1_1_NAND2_NUM122_OUT), .A2 (XNOR_1_2_NAND2_NUM122_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM122 (.ZN (N504), .A1 (XNOR_1_3_NAND2_NUM122_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM123_OUT, XNOR_1_2_NAND2_NUM123_OUT, XNOR_1_3_NAND2_NUM123_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM123 (.ZN (XNOR_1_1_NAND2_NUM123_OUT), .A1 (N416), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM123 (.ZN (XNOR_1_2_NAND2_NUM123_OUT), .A1 (GND), .A2 (N417));
      NOR2_X1 XNOR_1_3_NAND2_NUM123 (.ZN (XNOR_1_3_NAND2_NUM123_OUT), .A1 (XNOR_1_1_NAND2_NUM123_OUT), .A2 (XNOR_1_2_NAND2_NUM123_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM123 (.ZN (N507), .A1 (XNOR_1_3_NAND2_NUM123_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM124_OUT, XNOR_1_2_NAND2_NUM124_OUT, XNOR_1_3_NAND2_NUM124_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM124 (.ZN (XNOR_1_1_NAND2_NUM124_OUT), .A1 (N418), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM124 (.ZN (XNOR_1_2_NAND2_NUM124_OUT), .A1 (GND), .A2 (N419));
      NOR2_X1 XNOR_1_3_NAND2_NUM124 (.ZN (XNOR_1_3_NAND2_NUM124_OUT), .A1 (XNOR_1_1_NAND2_NUM124_OUT), .A2 (XNOR_1_2_NAND2_NUM124_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM124 (.ZN (N510), .A1 (XNOR_1_3_NAND2_NUM124_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM125_OUT, XNOR_1_2_NAND2_NUM125_OUT, XNOR_1_3_NAND2_NUM125_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM125 (.ZN (XNOR_1_1_NAND2_NUM125_OUT), .A1 (N420), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM125 (.ZN (XNOR_1_2_NAND2_NUM125_OUT), .A1 (GND), .A2 (N421));
      NOR2_X1 XNOR_1_3_NAND2_NUM125 (.ZN (XNOR_1_3_NAND2_NUM125_OUT), .A1 (XNOR_1_1_NAND2_NUM125_OUT), .A2 (XNOR_1_2_NAND2_NUM125_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM125 (.ZN (N513), .A1 (XNOR_1_3_NAND2_NUM125_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM126_OUT, XNOR_1_2_NAND2_NUM126_OUT, XNOR_1_3_NAND2_NUM126_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM126 (.ZN (XNOR_1_1_NAND2_NUM126_OUT), .A1 (N422), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM126 (.ZN (XNOR_1_2_NAND2_NUM126_OUT), .A1 (GND), .A2 (N423));
      NOR2_X1 XNOR_1_3_NAND2_NUM126 (.ZN (XNOR_1_3_NAND2_NUM126_OUT), .A1 (XNOR_1_1_NAND2_NUM126_OUT), .A2 (XNOR_1_2_NAND2_NUM126_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM126 (.ZN (N516), .A1 (XNOR_1_3_NAND2_NUM126_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM127_OUT, XNOR_1_2_NAND2_NUM127_OUT, XNOR_1_3_NAND2_NUM127_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM127 (.ZN (XNOR_1_1_NAND2_NUM127_OUT), .A1 (N424), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM127 (.ZN (XNOR_1_2_NAND2_NUM127_OUT), .A1 (GND), .A2 (N425));
      NOR2_X1 XNOR_1_3_NAND2_NUM127 (.ZN (XNOR_1_3_NAND2_NUM127_OUT), .A1 (XNOR_1_1_NAND2_NUM127_OUT), .A2 (XNOR_1_2_NAND2_NUM127_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM127 (.ZN (N519), .A1 (XNOR_1_3_NAND2_NUM127_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM128_OUT, XNOR_1_2_NAND2_NUM128_OUT, XNOR_1_3_NAND2_NUM128_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM128 (.ZN (XNOR_1_1_NAND2_NUM128_OUT), .A1 (N426), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM128 (.ZN (XNOR_1_2_NAND2_NUM128_OUT), .A1 (GND), .A2 (N429));
      NOR2_X1 XNOR_1_3_NAND2_NUM128 (.ZN (XNOR_1_3_NAND2_NUM128_OUT), .A1 (XNOR_1_1_NAND2_NUM128_OUT), .A2 (XNOR_1_2_NAND2_NUM128_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM128 (.ZN (N522), .A1 (XNOR_1_3_NAND2_NUM128_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM129_OUT, XNOR_1_2_NAND2_NUM129_OUT, XNOR_1_3_NAND2_NUM129_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM129 (.ZN (XNOR_1_1_NAND2_NUM129_OUT), .A1 (N432), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM129 (.ZN (XNOR_1_2_NAND2_NUM129_OUT), .A1 (GND), .A2 (N435));
      NOR2_X1 XNOR_1_3_NAND2_NUM129 (.ZN (XNOR_1_3_NAND2_NUM129_OUT), .A1 (XNOR_1_1_NAND2_NUM129_OUT), .A2 (XNOR_1_2_NAND2_NUM129_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM129 (.ZN (N525), .A1 (XNOR_1_3_NAND2_NUM129_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM130_OUT, XNOR_1_2_NAND2_NUM130_OUT, XNOR_1_3_NAND2_NUM130_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM130 (.ZN (XNOR_1_1_NAND2_NUM130_OUT), .A1 (N438), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM130 (.ZN (XNOR_1_2_NAND2_NUM130_OUT), .A1 (GND), .A2 (N441));
      NOR2_X1 XNOR_1_3_NAND2_NUM130 (.ZN (XNOR_1_3_NAND2_NUM130_OUT), .A1 (XNOR_1_1_NAND2_NUM130_OUT), .A2 (XNOR_1_2_NAND2_NUM130_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM130 (.ZN (N528), .A1 (XNOR_1_3_NAND2_NUM130_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM131_OUT, XNOR_1_2_NAND2_NUM131_OUT, XNOR_1_3_NAND2_NUM131_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM131 (.ZN (XNOR_1_1_NAND2_NUM131_OUT), .A1 (N444), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM131 (.ZN (XNOR_1_2_NAND2_NUM131_OUT), .A1 (GND), .A2 (N447));
      NOR2_X1 XNOR_1_3_NAND2_NUM131 (.ZN (XNOR_1_3_NAND2_NUM131_OUT), .A1 (XNOR_1_1_NAND2_NUM131_OUT), .A2 (XNOR_1_2_NAND2_NUM131_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM131 (.ZN (N531), .A1 (XNOR_1_3_NAND2_NUM131_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM132_OUT, XNOR_1_2_NAND2_NUM132_OUT, XNOR_1_3_NAND2_NUM132_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM132 (.ZN (XNOR_1_1_NAND2_NUM132_OUT), .A1 (N450), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM132 (.ZN (XNOR_1_2_NAND2_NUM132_OUT), .A1 (GND), .A2 (N453));
      NOR2_X1 XNOR_1_3_NAND2_NUM132 (.ZN (XNOR_1_3_NAND2_NUM132_OUT), .A1 (XNOR_1_1_NAND2_NUM132_OUT), .A2 (XNOR_1_2_NAND2_NUM132_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM132 (.ZN (N534), .A1 (XNOR_1_3_NAND2_NUM132_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM133_OUT, XNOR_1_2_NAND2_NUM133_OUT, XNOR_1_3_NAND2_NUM133_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM133 (.ZN (XNOR_1_1_NAND2_NUM133_OUT), .A1 (N456), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM133 (.ZN (XNOR_1_2_NAND2_NUM133_OUT), .A1 (GND), .A2 (N459));
      NOR2_X1 XNOR_1_3_NAND2_NUM133 (.ZN (XNOR_1_3_NAND2_NUM133_OUT), .A1 (XNOR_1_1_NAND2_NUM133_OUT), .A2 (XNOR_1_2_NAND2_NUM133_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM133 (.ZN (N537), .A1 (XNOR_1_3_NAND2_NUM133_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM134_OUT, XNOR_1_2_NAND2_NUM134_OUT, XNOR_1_3_NAND2_NUM134_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM134 (.ZN (XNOR_1_1_NAND2_NUM134_OUT), .A1 (N462), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM134 (.ZN (XNOR_1_2_NAND2_NUM134_OUT), .A1 (GND), .A2 (N465));
      NOR2_X1 XNOR_1_3_NAND2_NUM134 (.ZN (XNOR_1_3_NAND2_NUM134_OUT), .A1 (XNOR_1_1_NAND2_NUM134_OUT), .A2 (XNOR_1_2_NAND2_NUM134_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM134 (.ZN (N540), .A1 (XNOR_1_3_NAND2_NUM134_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM135_OUT, XNOR_1_2_NAND2_NUM135_OUT, XNOR_1_3_NAND2_NUM135_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM135 (.ZN (XNOR_1_1_NAND2_NUM135_OUT), .A1 (N468), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM135 (.ZN (XNOR_1_2_NAND2_NUM135_OUT), .A1 (GND), .A2 (N471));
      NOR2_X1 XNOR_1_3_NAND2_NUM135 (.ZN (XNOR_1_3_NAND2_NUM135_OUT), .A1 (XNOR_1_1_NAND2_NUM135_OUT), .A2 (XNOR_1_2_NAND2_NUM135_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM135 (.ZN (N543), .A1 (XNOR_1_3_NAND2_NUM135_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM136_OUT, XNOR_1_2_NAND2_NUM136_OUT, XNOR_1_3_NAND2_NUM136_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM136 (.ZN (XNOR_1_1_NAND2_NUM136_OUT), .A1 (N474), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM136 (.ZN (XNOR_1_2_NAND2_NUM136_OUT), .A1 (GND), .A2 (N477));
      NOR2_X1 XNOR_1_3_NAND2_NUM136 (.ZN (XNOR_1_3_NAND2_NUM136_OUT), .A1 (XNOR_1_1_NAND2_NUM136_OUT), .A2 (XNOR_1_2_NAND2_NUM136_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM136 (.ZN (N546), .A1 (XNOR_1_3_NAND2_NUM136_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM137_OUT, XNOR_1_2_NAND2_NUM137_OUT, XNOR_1_3_NAND2_NUM137_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM137 (.ZN (XNOR_1_1_NAND2_NUM137_OUT), .A1 (N480), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM137 (.ZN (XNOR_1_2_NAND2_NUM137_OUT), .A1 (GND), .A2 (N483));
      NOR2_X1 XNOR_1_3_NAND2_NUM137 (.ZN (XNOR_1_3_NAND2_NUM137_OUT), .A1 (XNOR_1_1_NAND2_NUM137_OUT), .A2 (XNOR_1_2_NAND2_NUM137_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM137 (.ZN (N549), .A1 (XNOR_1_3_NAND2_NUM137_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM138_OUT, XNOR_1_2_NAND2_NUM138_OUT, XNOR_1_3_NAND2_NUM138_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM138 (.ZN (XNOR_1_1_NAND2_NUM138_OUT), .A1 (N486), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM138 (.ZN (XNOR_1_2_NAND2_NUM138_OUT), .A1 (GND), .A2 (N489));
      NOR2_X1 XNOR_1_3_NAND2_NUM138 (.ZN (XNOR_1_3_NAND2_NUM138_OUT), .A1 (XNOR_1_1_NAND2_NUM138_OUT), .A2 (XNOR_1_2_NAND2_NUM138_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM138 (.ZN (N552), .A1 (XNOR_1_3_NAND2_NUM138_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM139_OUT, XNOR_1_2_NAND2_NUM139_OUT, XNOR_1_3_NAND2_NUM139_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM139 (.ZN (XNOR_1_1_NAND2_NUM139_OUT), .A1 (N492), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM139 (.ZN (XNOR_1_2_NAND2_NUM139_OUT), .A1 (GND), .A2 (N495));
      NOR2_X1 XNOR_1_3_NAND2_NUM139 (.ZN (XNOR_1_3_NAND2_NUM139_OUT), .A1 (XNOR_1_1_NAND2_NUM139_OUT), .A2 (XNOR_1_2_NAND2_NUM139_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM139 (.ZN (N555), .A1 (XNOR_1_3_NAND2_NUM139_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM140_OUT, XNOR_1_2_NAND2_NUM140_OUT, XNOR_1_3_NAND2_NUM140_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM140 (.ZN (XNOR_1_1_NAND2_NUM140_OUT), .A1 (N498), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM140 (.ZN (XNOR_1_2_NAND2_NUM140_OUT), .A1 (GND), .A2 (N501));
      NOR2_X1 XNOR_1_3_NAND2_NUM140 (.ZN (XNOR_1_3_NAND2_NUM140_OUT), .A1 (XNOR_1_1_NAND2_NUM140_OUT), .A2 (XNOR_1_2_NAND2_NUM140_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM140 (.ZN (N558), .A1 (XNOR_1_3_NAND2_NUM140_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM141_OUT, XNOR_1_2_NAND2_NUM141_OUT, XNOR_1_3_NAND2_NUM141_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM141 (.ZN (XNOR_1_1_NAND2_NUM141_OUT), .A1 (N504), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM141 (.ZN (XNOR_1_2_NAND2_NUM141_OUT), .A1 (GND), .A2 (N507));
      NOR2_X1 XNOR_1_3_NAND2_NUM141 (.ZN (XNOR_1_3_NAND2_NUM141_OUT), .A1 (XNOR_1_1_NAND2_NUM141_OUT), .A2 (XNOR_1_2_NAND2_NUM141_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM141 (.ZN (N561), .A1 (XNOR_1_3_NAND2_NUM141_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM142_OUT, XNOR_1_2_NAND2_NUM142_OUT, XNOR_1_3_NAND2_NUM142_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM142 (.ZN (XNOR_1_1_NAND2_NUM142_OUT), .A1 (N510), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM142 (.ZN (XNOR_1_2_NAND2_NUM142_OUT), .A1 (GND), .A2 (N513));
      NOR2_X1 XNOR_1_3_NAND2_NUM142 (.ZN (XNOR_1_3_NAND2_NUM142_OUT), .A1 (XNOR_1_1_NAND2_NUM142_OUT), .A2 (XNOR_1_2_NAND2_NUM142_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM142 (.ZN (N564), .A1 (XNOR_1_3_NAND2_NUM142_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM143_OUT, XNOR_1_2_NAND2_NUM143_OUT, XNOR_1_3_NAND2_NUM143_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM143 (.ZN (XNOR_1_1_NAND2_NUM143_OUT), .A1 (N516), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM143 (.ZN (XNOR_1_2_NAND2_NUM143_OUT), .A1 (GND), .A2 (N519));
      NOR2_X1 XNOR_1_3_NAND2_NUM143 (.ZN (XNOR_1_3_NAND2_NUM143_OUT), .A1 (XNOR_1_1_NAND2_NUM143_OUT), .A2 (XNOR_1_2_NAND2_NUM143_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM143 (.ZN (N567), .A1 (XNOR_1_3_NAND2_NUM143_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM144_OUT, XNOR_1_2_NAND2_NUM144_OUT, XNOR_1_3_NAND2_NUM144_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM144 (.ZN (XNOR_1_1_NAND2_NUM144_OUT), .A1 (N426), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM144 (.ZN (XNOR_1_2_NAND2_NUM144_OUT), .A1 (GND), .A2 (N522));
      NOR2_X1 XNOR_1_3_NAND2_NUM144 (.ZN (XNOR_1_3_NAND2_NUM144_OUT), .A1 (XNOR_1_1_NAND2_NUM144_OUT), .A2 (XNOR_1_2_NAND2_NUM144_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM144 (.ZN (N570), .A1 (XNOR_1_3_NAND2_NUM144_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM145_OUT, XNOR_1_2_NAND2_NUM145_OUT, XNOR_1_3_NAND2_NUM145_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM145 (.ZN (XNOR_1_1_NAND2_NUM145_OUT), .A1 (N429), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM145 (.ZN (XNOR_1_2_NAND2_NUM145_OUT), .A1 (GND), .A2 (N522));
      NOR2_X1 XNOR_1_3_NAND2_NUM145 (.ZN (XNOR_1_3_NAND2_NUM145_OUT), .A1 (XNOR_1_1_NAND2_NUM145_OUT), .A2 (XNOR_1_2_NAND2_NUM145_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM145 (.ZN (N571), .A1 (XNOR_1_3_NAND2_NUM145_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM146_OUT, XNOR_1_2_NAND2_NUM146_OUT, XNOR_1_3_NAND2_NUM146_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM146 (.ZN (XNOR_1_1_NAND2_NUM146_OUT), .A1 (N432), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM146 (.ZN (XNOR_1_2_NAND2_NUM146_OUT), .A1 (GND), .A2 (N525));
      NOR2_X1 XNOR_1_3_NAND2_NUM146 (.ZN (XNOR_1_3_NAND2_NUM146_OUT), .A1 (XNOR_1_1_NAND2_NUM146_OUT), .A2 (XNOR_1_2_NAND2_NUM146_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM146 (.ZN (N572), .A1 (XNOR_1_3_NAND2_NUM146_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM147_OUT, XNOR_1_2_NAND2_NUM147_OUT, XNOR_1_3_NAND2_NUM147_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM147 (.ZN (XNOR_1_1_NAND2_NUM147_OUT), .A1 (N435), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM147 (.ZN (XNOR_1_2_NAND2_NUM147_OUT), .A1 (GND), .A2 (N525));
      NOR2_X1 XNOR_1_3_NAND2_NUM147 (.ZN (XNOR_1_3_NAND2_NUM147_OUT), .A1 (XNOR_1_1_NAND2_NUM147_OUT), .A2 (XNOR_1_2_NAND2_NUM147_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM147 (.ZN (N573), .A1 (XNOR_1_3_NAND2_NUM147_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM148_OUT, XNOR_1_2_NAND2_NUM148_OUT, XNOR_1_3_NAND2_NUM148_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM148 (.ZN (XNOR_1_1_NAND2_NUM148_OUT), .A1 (N438), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM148 (.ZN (XNOR_1_2_NAND2_NUM148_OUT), .A1 (GND), .A2 (N528));
      NOR2_X1 XNOR_1_3_NAND2_NUM148 (.ZN (XNOR_1_3_NAND2_NUM148_OUT), .A1 (XNOR_1_1_NAND2_NUM148_OUT), .A2 (XNOR_1_2_NAND2_NUM148_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM148 (.ZN (N574), .A1 (XNOR_1_3_NAND2_NUM148_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM149_OUT, XNOR_1_2_NAND2_NUM149_OUT, XNOR_1_3_NAND2_NUM149_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM149 (.ZN (XNOR_1_1_NAND2_NUM149_OUT), .A1 (N441), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM149 (.ZN (XNOR_1_2_NAND2_NUM149_OUT), .A1 (GND), .A2 (N528));
      NOR2_X1 XNOR_1_3_NAND2_NUM149 (.ZN (XNOR_1_3_NAND2_NUM149_OUT), .A1 (XNOR_1_1_NAND2_NUM149_OUT), .A2 (XNOR_1_2_NAND2_NUM149_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM149 (.ZN (N575), .A1 (XNOR_1_3_NAND2_NUM149_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM150_OUT, XNOR_1_2_NAND2_NUM150_OUT, XNOR_1_3_NAND2_NUM150_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM150 (.ZN (XNOR_1_1_NAND2_NUM150_OUT), .A1 (N444), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM150 (.ZN (XNOR_1_2_NAND2_NUM150_OUT), .A1 (GND), .A2 (N531));
      NOR2_X1 XNOR_1_3_NAND2_NUM150 (.ZN (XNOR_1_3_NAND2_NUM150_OUT), .A1 (XNOR_1_1_NAND2_NUM150_OUT), .A2 (XNOR_1_2_NAND2_NUM150_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM150 (.ZN (N576), .A1 (XNOR_1_3_NAND2_NUM150_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM151_OUT, XNOR_1_2_NAND2_NUM151_OUT, XNOR_1_3_NAND2_NUM151_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM151 (.ZN (XNOR_1_1_NAND2_NUM151_OUT), .A1 (N447), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM151 (.ZN (XNOR_1_2_NAND2_NUM151_OUT), .A1 (GND), .A2 (N531));
      NOR2_X1 XNOR_1_3_NAND2_NUM151 (.ZN (XNOR_1_3_NAND2_NUM151_OUT), .A1 (XNOR_1_1_NAND2_NUM151_OUT), .A2 (XNOR_1_2_NAND2_NUM151_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM151 (.ZN (N577), .A1 (XNOR_1_3_NAND2_NUM151_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM152_OUT, XNOR_1_2_NAND2_NUM152_OUT, XNOR_1_3_NAND2_NUM152_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM152 (.ZN (XNOR_1_1_NAND2_NUM152_OUT), .A1 (N450), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM152 (.ZN (XNOR_1_2_NAND2_NUM152_OUT), .A1 (GND), .A2 (N534));
      NOR2_X1 XNOR_1_3_NAND2_NUM152 (.ZN (XNOR_1_3_NAND2_NUM152_OUT), .A1 (XNOR_1_1_NAND2_NUM152_OUT), .A2 (XNOR_1_2_NAND2_NUM152_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM152 (.ZN (N578), .A1 (XNOR_1_3_NAND2_NUM152_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM153_OUT, XNOR_1_2_NAND2_NUM153_OUT, XNOR_1_3_NAND2_NUM153_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM153 (.ZN (XNOR_1_1_NAND2_NUM153_OUT), .A1 (N453), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM153 (.ZN (XNOR_1_2_NAND2_NUM153_OUT), .A1 (GND), .A2 (N534));
      NOR2_X1 XNOR_1_3_NAND2_NUM153 (.ZN (XNOR_1_3_NAND2_NUM153_OUT), .A1 (XNOR_1_1_NAND2_NUM153_OUT), .A2 (XNOR_1_2_NAND2_NUM153_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM153 (.ZN (N579), .A1 (XNOR_1_3_NAND2_NUM153_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM154_OUT, XNOR_1_2_NAND2_NUM154_OUT, XNOR_1_3_NAND2_NUM154_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM154 (.ZN (XNOR_1_1_NAND2_NUM154_OUT), .A1 (N456), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM154 (.ZN (XNOR_1_2_NAND2_NUM154_OUT), .A1 (GND), .A2 (N537));
      NOR2_X1 XNOR_1_3_NAND2_NUM154 (.ZN (XNOR_1_3_NAND2_NUM154_OUT), .A1 (XNOR_1_1_NAND2_NUM154_OUT), .A2 (XNOR_1_2_NAND2_NUM154_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM154 (.ZN (N580), .A1 (XNOR_1_3_NAND2_NUM154_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM155_OUT, XNOR_1_2_NAND2_NUM155_OUT, XNOR_1_3_NAND2_NUM155_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM155 (.ZN (XNOR_1_1_NAND2_NUM155_OUT), .A1 (N459), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM155 (.ZN (XNOR_1_2_NAND2_NUM155_OUT), .A1 (GND), .A2 (N537));
      NOR2_X1 XNOR_1_3_NAND2_NUM155 (.ZN (XNOR_1_3_NAND2_NUM155_OUT), .A1 (XNOR_1_1_NAND2_NUM155_OUT), .A2 (XNOR_1_2_NAND2_NUM155_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM155 (.ZN (N581), .A1 (XNOR_1_3_NAND2_NUM155_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM156_OUT, XNOR_1_2_NAND2_NUM156_OUT, XNOR_1_3_NAND2_NUM156_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM156 (.ZN (XNOR_1_1_NAND2_NUM156_OUT), .A1 (N462), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM156 (.ZN (XNOR_1_2_NAND2_NUM156_OUT), .A1 (GND), .A2 (N540));
      NOR2_X1 XNOR_1_3_NAND2_NUM156 (.ZN (XNOR_1_3_NAND2_NUM156_OUT), .A1 (XNOR_1_1_NAND2_NUM156_OUT), .A2 (XNOR_1_2_NAND2_NUM156_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM156 (.ZN (N582), .A1 (XNOR_1_3_NAND2_NUM156_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM157_OUT, XNOR_1_2_NAND2_NUM157_OUT, XNOR_1_3_NAND2_NUM157_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM157 (.ZN (XNOR_1_1_NAND2_NUM157_OUT), .A1 (N465), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM157 (.ZN (XNOR_1_2_NAND2_NUM157_OUT), .A1 (GND), .A2 (N540));
      NOR2_X1 XNOR_1_3_NAND2_NUM157 (.ZN (XNOR_1_3_NAND2_NUM157_OUT), .A1 (XNOR_1_1_NAND2_NUM157_OUT), .A2 (XNOR_1_2_NAND2_NUM157_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM157 (.ZN (N583), .A1 (XNOR_1_3_NAND2_NUM157_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM158_OUT, XNOR_1_2_NAND2_NUM158_OUT, XNOR_1_3_NAND2_NUM158_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM158 (.ZN (XNOR_1_1_NAND2_NUM158_OUT), .A1 (N468), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM158 (.ZN (XNOR_1_2_NAND2_NUM158_OUT), .A1 (GND), .A2 (N543));
      NOR2_X1 XNOR_1_3_NAND2_NUM158 (.ZN (XNOR_1_3_NAND2_NUM158_OUT), .A1 (XNOR_1_1_NAND2_NUM158_OUT), .A2 (XNOR_1_2_NAND2_NUM158_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM158 (.ZN (N584), .A1 (XNOR_1_3_NAND2_NUM158_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM159_OUT, XNOR_1_2_NAND2_NUM159_OUT, XNOR_1_3_NAND2_NUM159_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM159 (.ZN (XNOR_1_1_NAND2_NUM159_OUT), .A1 (N471), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM159 (.ZN (XNOR_1_2_NAND2_NUM159_OUT), .A1 (GND), .A2 (N543));
      NOR2_X1 XNOR_1_3_NAND2_NUM159 (.ZN (XNOR_1_3_NAND2_NUM159_OUT), .A1 (XNOR_1_1_NAND2_NUM159_OUT), .A2 (XNOR_1_2_NAND2_NUM159_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM159 (.ZN (N585), .A1 (XNOR_1_3_NAND2_NUM159_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM160_OUT, XNOR_1_2_NAND2_NUM160_OUT, XNOR_1_3_NAND2_NUM160_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM160 (.ZN (XNOR_1_1_NAND2_NUM160_OUT), .A1 (N474), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM160 (.ZN (XNOR_1_2_NAND2_NUM160_OUT), .A1 (GND), .A2 (N546));
      NOR2_X1 XNOR_1_3_NAND2_NUM160 (.ZN (XNOR_1_3_NAND2_NUM160_OUT), .A1 (XNOR_1_1_NAND2_NUM160_OUT), .A2 (XNOR_1_2_NAND2_NUM160_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM160 (.ZN (N586), .A1 (XNOR_1_3_NAND2_NUM160_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM161_OUT, XNOR_1_2_NAND2_NUM161_OUT, XNOR_1_3_NAND2_NUM161_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM161 (.ZN (XNOR_1_1_NAND2_NUM161_OUT), .A1 (N477), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM161 (.ZN (XNOR_1_2_NAND2_NUM161_OUT), .A1 (GND), .A2 (N546));
      NOR2_X1 XNOR_1_3_NAND2_NUM161 (.ZN (XNOR_1_3_NAND2_NUM161_OUT), .A1 (XNOR_1_1_NAND2_NUM161_OUT), .A2 (XNOR_1_2_NAND2_NUM161_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM161 (.ZN (N587), .A1 (XNOR_1_3_NAND2_NUM161_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM162_OUT, XNOR_1_2_NAND2_NUM162_OUT, XNOR_1_3_NAND2_NUM162_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM162 (.ZN (XNOR_1_1_NAND2_NUM162_OUT), .A1 (N480), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM162 (.ZN (XNOR_1_2_NAND2_NUM162_OUT), .A1 (GND), .A2 (N549));
      NOR2_X1 XNOR_1_3_NAND2_NUM162 (.ZN (XNOR_1_3_NAND2_NUM162_OUT), .A1 (XNOR_1_1_NAND2_NUM162_OUT), .A2 (XNOR_1_2_NAND2_NUM162_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM162 (.ZN (N588), .A1 (XNOR_1_3_NAND2_NUM162_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM163_OUT, XNOR_1_2_NAND2_NUM163_OUT, XNOR_1_3_NAND2_NUM163_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM163 (.ZN (XNOR_1_1_NAND2_NUM163_OUT), .A1 (N483), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM163 (.ZN (XNOR_1_2_NAND2_NUM163_OUT), .A1 (GND), .A2 (N549));
      NOR2_X1 XNOR_1_3_NAND2_NUM163 (.ZN (XNOR_1_3_NAND2_NUM163_OUT), .A1 (XNOR_1_1_NAND2_NUM163_OUT), .A2 (XNOR_1_2_NAND2_NUM163_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM163 (.ZN (N589), .A1 (XNOR_1_3_NAND2_NUM163_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM164_OUT, XNOR_1_2_NAND2_NUM164_OUT, XNOR_1_3_NAND2_NUM164_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM164 (.ZN (XNOR_1_1_NAND2_NUM164_OUT), .A1 (N486), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM164 (.ZN (XNOR_1_2_NAND2_NUM164_OUT), .A1 (GND), .A2 (N552));
      NOR2_X1 XNOR_1_3_NAND2_NUM164 (.ZN (XNOR_1_3_NAND2_NUM164_OUT), .A1 (XNOR_1_1_NAND2_NUM164_OUT), .A2 (XNOR_1_2_NAND2_NUM164_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM164 (.ZN (N590), .A1 (XNOR_1_3_NAND2_NUM164_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM165_OUT, XNOR_1_2_NAND2_NUM165_OUT, XNOR_1_3_NAND2_NUM165_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM165 (.ZN (XNOR_1_1_NAND2_NUM165_OUT), .A1 (N489), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM165 (.ZN (XNOR_1_2_NAND2_NUM165_OUT), .A1 (GND), .A2 (N552));
      NOR2_X1 XNOR_1_3_NAND2_NUM165 (.ZN (XNOR_1_3_NAND2_NUM165_OUT), .A1 (XNOR_1_1_NAND2_NUM165_OUT), .A2 (XNOR_1_2_NAND2_NUM165_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM165 (.ZN (N591), .A1 (XNOR_1_3_NAND2_NUM165_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM166_OUT, XNOR_1_2_NAND2_NUM166_OUT, XNOR_1_3_NAND2_NUM166_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM166 (.ZN (XNOR_1_1_NAND2_NUM166_OUT), .A1 (N492), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM166 (.ZN (XNOR_1_2_NAND2_NUM166_OUT), .A1 (GND), .A2 (N555));
      NOR2_X1 XNOR_1_3_NAND2_NUM166 (.ZN (XNOR_1_3_NAND2_NUM166_OUT), .A1 (XNOR_1_1_NAND2_NUM166_OUT), .A2 (XNOR_1_2_NAND2_NUM166_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM166 (.ZN (N592), .A1 (XNOR_1_3_NAND2_NUM166_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM167_OUT, XNOR_1_2_NAND2_NUM167_OUT, XNOR_1_3_NAND2_NUM167_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM167 (.ZN (XNOR_1_1_NAND2_NUM167_OUT), .A1 (N495), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM167 (.ZN (XNOR_1_2_NAND2_NUM167_OUT), .A1 (GND), .A2 (N555));
      NOR2_X1 XNOR_1_3_NAND2_NUM167 (.ZN (XNOR_1_3_NAND2_NUM167_OUT), .A1 (XNOR_1_1_NAND2_NUM167_OUT), .A2 (XNOR_1_2_NAND2_NUM167_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM167 (.ZN (N593), .A1 (XNOR_1_3_NAND2_NUM167_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM168_OUT, XNOR_1_2_NAND2_NUM168_OUT, XNOR_1_3_NAND2_NUM168_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM168 (.ZN (XNOR_1_1_NAND2_NUM168_OUT), .A1 (N498), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM168 (.ZN (XNOR_1_2_NAND2_NUM168_OUT), .A1 (GND), .A2 (N558));
      NOR2_X1 XNOR_1_3_NAND2_NUM168 (.ZN (XNOR_1_3_NAND2_NUM168_OUT), .A1 (XNOR_1_1_NAND2_NUM168_OUT), .A2 (XNOR_1_2_NAND2_NUM168_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM168 (.ZN (N594), .A1 (XNOR_1_3_NAND2_NUM168_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM169_OUT, XNOR_1_2_NAND2_NUM169_OUT, XNOR_1_3_NAND2_NUM169_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM169 (.ZN (XNOR_1_1_NAND2_NUM169_OUT), .A1 (N501), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM169 (.ZN (XNOR_1_2_NAND2_NUM169_OUT), .A1 (GND), .A2 (N558));
      NOR2_X1 XNOR_1_3_NAND2_NUM169 (.ZN (XNOR_1_3_NAND2_NUM169_OUT), .A1 (XNOR_1_1_NAND2_NUM169_OUT), .A2 (XNOR_1_2_NAND2_NUM169_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM169 (.ZN (N595), .A1 (XNOR_1_3_NAND2_NUM169_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM170_OUT, XNOR_1_2_NAND2_NUM170_OUT, XNOR_1_3_NAND2_NUM170_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM170 (.ZN (XNOR_1_1_NAND2_NUM170_OUT), .A1 (N504), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM170 (.ZN (XNOR_1_2_NAND2_NUM170_OUT), .A1 (GND), .A2 (N561));
      NOR2_X1 XNOR_1_3_NAND2_NUM170 (.ZN (XNOR_1_3_NAND2_NUM170_OUT), .A1 (XNOR_1_1_NAND2_NUM170_OUT), .A2 (XNOR_1_2_NAND2_NUM170_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM170 (.ZN (N596), .A1 (XNOR_1_3_NAND2_NUM170_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM171_OUT, XNOR_1_2_NAND2_NUM171_OUT, XNOR_1_3_NAND2_NUM171_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM171 (.ZN (XNOR_1_1_NAND2_NUM171_OUT), .A1 (N507), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM171 (.ZN (XNOR_1_2_NAND2_NUM171_OUT), .A1 (GND), .A2 (N561));
      NOR2_X1 XNOR_1_3_NAND2_NUM171 (.ZN (XNOR_1_3_NAND2_NUM171_OUT), .A1 (XNOR_1_1_NAND2_NUM171_OUT), .A2 (XNOR_1_2_NAND2_NUM171_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM171 (.ZN (N597), .A1 (XNOR_1_3_NAND2_NUM171_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM172_OUT, XNOR_1_2_NAND2_NUM172_OUT, XNOR_1_3_NAND2_NUM172_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM172 (.ZN (XNOR_1_1_NAND2_NUM172_OUT), .A1 (N510), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM172 (.ZN (XNOR_1_2_NAND2_NUM172_OUT), .A1 (GND), .A2 (N564));
      NOR2_X1 XNOR_1_3_NAND2_NUM172 (.ZN (XNOR_1_3_NAND2_NUM172_OUT), .A1 (XNOR_1_1_NAND2_NUM172_OUT), .A2 (XNOR_1_2_NAND2_NUM172_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM172 (.ZN (N598), .A1 (XNOR_1_3_NAND2_NUM172_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM173_OUT, XNOR_1_2_NAND2_NUM173_OUT, XNOR_1_3_NAND2_NUM173_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM173 (.ZN (XNOR_1_1_NAND2_NUM173_OUT), .A1 (N513), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM173 (.ZN (XNOR_1_2_NAND2_NUM173_OUT), .A1 (GND), .A2 (N564));
      NOR2_X1 XNOR_1_3_NAND2_NUM173 (.ZN (XNOR_1_3_NAND2_NUM173_OUT), .A1 (XNOR_1_1_NAND2_NUM173_OUT), .A2 (XNOR_1_2_NAND2_NUM173_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM173 (.ZN (N599), .A1 (XNOR_1_3_NAND2_NUM173_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM174_OUT, XNOR_1_2_NAND2_NUM174_OUT, XNOR_1_3_NAND2_NUM174_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM174 (.ZN (XNOR_1_1_NAND2_NUM174_OUT), .A1 (N516), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM174 (.ZN (XNOR_1_2_NAND2_NUM174_OUT), .A1 (GND), .A2 (N567));
      NOR2_X1 XNOR_1_3_NAND2_NUM174 (.ZN (XNOR_1_3_NAND2_NUM174_OUT), .A1 (XNOR_1_1_NAND2_NUM174_OUT), .A2 (XNOR_1_2_NAND2_NUM174_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM174 (.ZN (N600), .A1 (XNOR_1_3_NAND2_NUM174_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM175_OUT, XNOR_1_2_NAND2_NUM175_OUT, XNOR_1_3_NAND2_NUM175_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM175 (.ZN (XNOR_1_1_NAND2_NUM175_OUT), .A1 (N519), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM175 (.ZN (XNOR_1_2_NAND2_NUM175_OUT), .A1 (GND), .A2 (N567));
      NOR2_X1 XNOR_1_3_NAND2_NUM175 (.ZN (XNOR_1_3_NAND2_NUM175_OUT), .A1 (XNOR_1_1_NAND2_NUM175_OUT), .A2 (XNOR_1_2_NAND2_NUM175_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM175 (.ZN (N601), .A1 (XNOR_1_3_NAND2_NUM175_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM176_OUT, XNOR_1_2_NAND2_NUM176_OUT, XNOR_1_3_NAND2_NUM176_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM176 (.ZN (XNOR_1_1_NAND2_NUM176_OUT), .A1 (N570), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM176 (.ZN (XNOR_1_2_NAND2_NUM176_OUT), .A1 (GND), .A2 (N571));
      NOR2_X1 XNOR_1_3_NAND2_NUM176 (.ZN (XNOR_1_3_NAND2_NUM176_OUT), .A1 (XNOR_1_1_NAND2_NUM176_OUT), .A2 (XNOR_1_2_NAND2_NUM176_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM176 (.ZN (N602), .A1 (XNOR_1_3_NAND2_NUM176_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM177_OUT, XNOR_1_2_NAND2_NUM177_OUT, XNOR_1_3_NAND2_NUM177_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM177 (.ZN (XNOR_1_1_NAND2_NUM177_OUT), .A1 (N572), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM177 (.ZN (XNOR_1_2_NAND2_NUM177_OUT), .A1 (GND), .A2 (N573));
      NOR2_X1 XNOR_1_3_NAND2_NUM177 (.ZN (XNOR_1_3_NAND2_NUM177_OUT), .A1 (XNOR_1_1_NAND2_NUM177_OUT), .A2 (XNOR_1_2_NAND2_NUM177_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM177 (.ZN (N607), .A1 (XNOR_1_3_NAND2_NUM177_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM178_OUT, XNOR_1_2_NAND2_NUM178_OUT, XNOR_1_3_NAND2_NUM178_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM178 (.ZN (XNOR_1_1_NAND2_NUM178_OUT), .A1 (N574), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM178 (.ZN (XNOR_1_2_NAND2_NUM178_OUT), .A1 (GND), .A2 (N575));
      NOR2_X1 XNOR_1_3_NAND2_NUM178 (.ZN (XNOR_1_3_NAND2_NUM178_OUT), .A1 (XNOR_1_1_NAND2_NUM178_OUT), .A2 (XNOR_1_2_NAND2_NUM178_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM178 (.ZN (N612), .A1 (XNOR_1_3_NAND2_NUM178_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM179_OUT, XNOR_1_2_NAND2_NUM179_OUT, XNOR_1_3_NAND2_NUM179_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM179 (.ZN (XNOR_1_1_NAND2_NUM179_OUT), .A1 (N576), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM179 (.ZN (XNOR_1_2_NAND2_NUM179_OUT), .A1 (GND), .A2 (N577));
      NOR2_X1 XNOR_1_3_NAND2_NUM179 (.ZN (XNOR_1_3_NAND2_NUM179_OUT), .A1 (XNOR_1_1_NAND2_NUM179_OUT), .A2 (XNOR_1_2_NAND2_NUM179_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM179 (.ZN (N617), .A1 (XNOR_1_3_NAND2_NUM179_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM180_OUT, XNOR_1_2_NAND2_NUM180_OUT, XNOR_1_3_NAND2_NUM180_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM180 (.ZN (XNOR_1_1_NAND2_NUM180_OUT), .A1 (N578), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM180 (.ZN (XNOR_1_2_NAND2_NUM180_OUT), .A1 (GND), .A2 (N579));
      NOR2_X1 XNOR_1_3_NAND2_NUM180 (.ZN (XNOR_1_3_NAND2_NUM180_OUT), .A1 (XNOR_1_1_NAND2_NUM180_OUT), .A2 (XNOR_1_2_NAND2_NUM180_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM180 (.ZN (N622), .A1 (XNOR_1_3_NAND2_NUM180_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM181_OUT, XNOR_1_2_NAND2_NUM181_OUT, XNOR_1_3_NAND2_NUM181_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM181 (.ZN (XNOR_1_1_NAND2_NUM181_OUT), .A1 (N580), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM181 (.ZN (XNOR_1_2_NAND2_NUM181_OUT), .A1 (GND), .A2 (N581));
      NOR2_X1 XNOR_1_3_NAND2_NUM181 (.ZN (XNOR_1_3_NAND2_NUM181_OUT), .A1 (XNOR_1_1_NAND2_NUM181_OUT), .A2 (XNOR_1_2_NAND2_NUM181_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM181 (.ZN (N627), .A1 (XNOR_1_3_NAND2_NUM181_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM182_OUT, XNOR_1_2_NAND2_NUM182_OUT, XNOR_1_3_NAND2_NUM182_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM182 (.ZN (XNOR_1_1_NAND2_NUM182_OUT), .A1 (N582), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM182 (.ZN (XNOR_1_2_NAND2_NUM182_OUT), .A1 (GND), .A2 (N583));
      NOR2_X1 XNOR_1_3_NAND2_NUM182 (.ZN (XNOR_1_3_NAND2_NUM182_OUT), .A1 (XNOR_1_1_NAND2_NUM182_OUT), .A2 (XNOR_1_2_NAND2_NUM182_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM182 (.ZN (N632), .A1 (XNOR_1_3_NAND2_NUM182_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM183_OUT, XNOR_1_2_NAND2_NUM183_OUT, XNOR_1_3_NAND2_NUM183_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM183 (.ZN (XNOR_1_1_NAND2_NUM183_OUT), .A1 (N584), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM183 (.ZN (XNOR_1_2_NAND2_NUM183_OUT), .A1 (GND), .A2 (N585));
      NOR2_X1 XNOR_1_3_NAND2_NUM183 (.ZN (XNOR_1_3_NAND2_NUM183_OUT), .A1 (XNOR_1_1_NAND2_NUM183_OUT), .A2 (XNOR_1_2_NAND2_NUM183_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM183 (.ZN (N637), .A1 (XNOR_1_3_NAND2_NUM183_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM184_OUT, XNOR_1_2_NAND2_NUM184_OUT, XNOR_1_3_NAND2_NUM184_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM184 (.ZN (XNOR_1_1_NAND2_NUM184_OUT), .A1 (N586), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM184 (.ZN (XNOR_1_2_NAND2_NUM184_OUT), .A1 (GND), .A2 (N587));
      NOR2_X1 XNOR_1_3_NAND2_NUM184 (.ZN (XNOR_1_3_NAND2_NUM184_OUT), .A1 (XNOR_1_1_NAND2_NUM184_OUT), .A2 (XNOR_1_2_NAND2_NUM184_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM184 (.ZN (N642), .A1 (XNOR_1_3_NAND2_NUM184_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM185_OUT, XNOR_1_2_NAND2_NUM185_OUT, XNOR_1_3_NAND2_NUM185_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM185 (.ZN (XNOR_1_1_NAND2_NUM185_OUT), .A1 (N588), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM185 (.ZN (XNOR_1_2_NAND2_NUM185_OUT), .A1 (GND), .A2 (N589));
      NOR2_X1 XNOR_1_3_NAND2_NUM185 (.ZN (XNOR_1_3_NAND2_NUM185_OUT), .A1 (XNOR_1_1_NAND2_NUM185_OUT), .A2 (XNOR_1_2_NAND2_NUM185_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM185 (.ZN (N645), .A1 (XNOR_1_3_NAND2_NUM185_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM186_OUT, XNOR_1_2_NAND2_NUM186_OUT, XNOR_1_3_NAND2_NUM186_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM186 (.ZN (XNOR_1_1_NAND2_NUM186_OUT), .A1 (N590), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM186 (.ZN (XNOR_1_2_NAND2_NUM186_OUT), .A1 (GND), .A2 (N591));
      NOR2_X1 XNOR_1_3_NAND2_NUM186 (.ZN (XNOR_1_3_NAND2_NUM186_OUT), .A1 (XNOR_1_1_NAND2_NUM186_OUT), .A2 (XNOR_1_2_NAND2_NUM186_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM186 (.ZN (N648), .A1 (XNOR_1_3_NAND2_NUM186_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM187_OUT, XNOR_1_2_NAND2_NUM187_OUT, XNOR_1_3_NAND2_NUM187_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM187 (.ZN (XNOR_1_1_NAND2_NUM187_OUT), .A1 (N592), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM187 (.ZN (XNOR_1_2_NAND2_NUM187_OUT), .A1 (GND), .A2 (N593));
      NOR2_X1 XNOR_1_3_NAND2_NUM187 (.ZN (XNOR_1_3_NAND2_NUM187_OUT), .A1 (XNOR_1_1_NAND2_NUM187_OUT), .A2 (XNOR_1_2_NAND2_NUM187_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM187 (.ZN (N651), .A1 (XNOR_1_3_NAND2_NUM187_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM188_OUT, XNOR_1_2_NAND2_NUM188_OUT, XNOR_1_3_NAND2_NUM188_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM188 (.ZN (XNOR_1_1_NAND2_NUM188_OUT), .A1 (N594), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM188 (.ZN (XNOR_1_2_NAND2_NUM188_OUT), .A1 (GND), .A2 (N595));
      NOR2_X1 XNOR_1_3_NAND2_NUM188 (.ZN (XNOR_1_3_NAND2_NUM188_OUT), .A1 (XNOR_1_1_NAND2_NUM188_OUT), .A2 (XNOR_1_2_NAND2_NUM188_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM188 (.ZN (N654), .A1 (XNOR_1_3_NAND2_NUM188_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM189_OUT, XNOR_1_2_NAND2_NUM189_OUT, XNOR_1_3_NAND2_NUM189_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM189 (.ZN (XNOR_1_1_NAND2_NUM189_OUT), .A1 (N596), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM189 (.ZN (XNOR_1_2_NAND2_NUM189_OUT), .A1 (GND), .A2 (N597));
      NOR2_X1 XNOR_1_3_NAND2_NUM189 (.ZN (XNOR_1_3_NAND2_NUM189_OUT), .A1 (XNOR_1_1_NAND2_NUM189_OUT), .A2 (XNOR_1_2_NAND2_NUM189_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM189 (.ZN (N657), .A1 (XNOR_1_3_NAND2_NUM189_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM190_OUT, XNOR_1_2_NAND2_NUM190_OUT, XNOR_1_3_NAND2_NUM190_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM190 (.ZN (XNOR_1_1_NAND2_NUM190_OUT), .A1 (N598), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM190 (.ZN (XNOR_1_2_NAND2_NUM190_OUT), .A1 (GND), .A2 (N599));
      NOR2_X1 XNOR_1_3_NAND2_NUM190 (.ZN (XNOR_1_3_NAND2_NUM190_OUT), .A1 (XNOR_1_1_NAND2_NUM190_OUT), .A2 (XNOR_1_2_NAND2_NUM190_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM190 (.ZN (N660), .A1 (XNOR_1_3_NAND2_NUM190_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM191_OUT, XNOR_1_2_NAND2_NUM191_OUT, XNOR_1_3_NAND2_NUM191_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM191 (.ZN (XNOR_1_1_NAND2_NUM191_OUT), .A1 (N600), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM191 (.ZN (XNOR_1_2_NAND2_NUM191_OUT), .A1 (GND), .A2 (N601));
      NOR2_X1 XNOR_1_3_NAND2_NUM191 (.ZN (XNOR_1_3_NAND2_NUM191_OUT), .A1 (XNOR_1_1_NAND2_NUM191_OUT), .A2 (XNOR_1_2_NAND2_NUM191_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM191 (.ZN (N663), .A1 (XNOR_1_3_NAND2_NUM191_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM192_OUT, XNOR_1_2_NAND2_NUM192_OUT, XNOR_1_3_NAND2_NUM192_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM192 (.ZN (XNOR_1_1_NAND2_NUM192_OUT), .A1 (N602), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM192 (.ZN (XNOR_1_2_NAND2_NUM192_OUT), .A1 (GND), .A2 (N607));
      NOR2_X1 XNOR_1_3_NAND2_NUM192 (.ZN (XNOR_1_3_NAND2_NUM192_OUT), .A1 (XNOR_1_1_NAND2_NUM192_OUT), .A2 (XNOR_1_2_NAND2_NUM192_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM192 (.ZN (N666), .A1 (XNOR_1_3_NAND2_NUM192_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM193_OUT, XNOR_1_2_NAND2_NUM193_OUT, XNOR_1_3_NAND2_NUM193_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM193 (.ZN (XNOR_1_1_NAND2_NUM193_OUT), .A1 (N612), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM193 (.ZN (XNOR_1_2_NAND2_NUM193_OUT), .A1 (GND), .A2 (N617));
      NOR2_X1 XNOR_1_3_NAND2_NUM193 (.ZN (XNOR_1_3_NAND2_NUM193_OUT), .A1 (XNOR_1_1_NAND2_NUM193_OUT), .A2 (XNOR_1_2_NAND2_NUM193_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM193 (.ZN (N669), .A1 (XNOR_1_3_NAND2_NUM193_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM194_OUT, XNOR_1_2_NAND2_NUM194_OUT, XNOR_1_3_NAND2_NUM194_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM194 (.ZN (XNOR_1_1_NAND2_NUM194_OUT), .A1 (N602), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM194 (.ZN (XNOR_1_2_NAND2_NUM194_OUT), .A1 (GND), .A2 (N612));
      NOR2_X1 XNOR_1_3_NAND2_NUM194 (.ZN (XNOR_1_3_NAND2_NUM194_OUT), .A1 (XNOR_1_1_NAND2_NUM194_OUT), .A2 (XNOR_1_2_NAND2_NUM194_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM194 (.ZN (N672), .A1 (XNOR_1_3_NAND2_NUM194_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM195_OUT, XNOR_1_2_NAND2_NUM195_OUT, XNOR_1_3_NAND2_NUM195_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM195 (.ZN (XNOR_1_1_NAND2_NUM195_OUT), .A1 (N607), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM195 (.ZN (XNOR_1_2_NAND2_NUM195_OUT), .A1 (GND), .A2 (N617));
      NOR2_X1 XNOR_1_3_NAND2_NUM195 (.ZN (XNOR_1_3_NAND2_NUM195_OUT), .A1 (XNOR_1_1_NAND2_NUM195_OUT), .A2 (XNOR_1_2_NAND2_NUM195_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM195 (.ZN (N675), .A1 (XNOR_1_3_NAND2_NUM195_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM196_OUT, XNOR_1_2_NAND2_NUM196_OUT, XNOR_1_3_NAND2_NUM196_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM196 (.ZN (XNOR_1_1_NAND2_NUM196_OUT), .A1 (N622), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM196 (.ZN (XNOR_1_2_NAND2_NUM196_OUT), .A1 (GND), .A2 (N627));
      NOR2_X1 XNOR_1_3_NAND2_NUM196 (.ZN (XNOR_1_3_NAND2_NUM196_OUT), .A1 (XNOR_1_1_NAND2_NUM196_OUT), .A2 (XNOR_1_2_NAND2_NUM196_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM196 (.ZN (N678), .A1 (XNOR_1_3_NAND2_NUM196_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM197_OUT, XNOR_1_2_NAND2_NUM197_OUT, XNOR_1_3_NAND2_NUM197_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM197 (.ZN (XNOR_1_1_NAND2_NUM197_OUT), .A1 (N632), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM197 (.ZN (XNOR_1_2_NAND2_NUM197_OUT), .A1 (GND), .A2 (N637));
      NOR2_X1 XNOR_1_3_NAND2_NUM197 (.ZN (XNOR_1_3_NAND2_NUM197_OUT), .A1 (XNOR_1_1_NAND2_NUM197_OUT), .A2 (XNOR_1_2_NAND2_NUM197_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM197 (.ZN (N681), .A1 (XNOR_1_3_NAND2_NUM197_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM198_OUT, XNOR_1_2_NAND2_NUM198_OUT, XNOR_1_3_NAND2_NUM198_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM198 (.ZN (XNOR_1_1_NAND2_NUM198_OUT), .A1 (N622), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM198 (.ZN (XNOR_1_2_NAND2_NUM198_OUT), .A1 (GND), .A2 (N632));
      NOR2_X1 XNOR_1_3_NAND2_NUM198 (.ZN (XNOR_1_3_NAND2_NUM198_OUT), .A1 (XNOR_1_1_NAND2_NUM198_OUT), .A2 (XNOR_1_2_NAND2_NUM198_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM198 (.ZN (N684), .A1 (XNOR_1_3_NAND2_NUM198_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM199_OUT, XNOR_1_2_NAND2_NUM199_OUT, XNOR_1_3_NAND2_NUM199_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM199 (.ZN (XNOR_1_1_NAND2_NUM199_OUT), .A1 (N627), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM199 (.ZN (XNOR_1_2_NAND2_NUM199_OUT), .A1 (GND), .A2 (N637));
      NOR2_X1 XNOR_1_3_NAND2_NUM199 (.ZN (XNOR_1_3_NAND2_NUM199_OUT), .A1 (XNOR_1_1_NAND2_NUM199_OUT), .A2 (XNOR_1_2_NAND2_NUM199_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM199 (.ZN (N687), .A1 (XNOR_1_3_NAND2_NUM199_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM200_OUT, XNOR_1_2_NAND2_NUM200_OUT, XNOR_1_3_NAND2_NUM200_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM200 (.ZN (XNOR_1_1_NAND2_NUM200_OUT), .A1 (N602), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM200 (.ZN (XNOR_1_2_NAND2_NUM200_OUT), .A1 (GND), .A2 (N666));
      NOR2_X1 XNOR_1_3_NAND2_NUM200 (.ZN (XNOR_1_3_NAND2_NUM200_OUT), .A1 (XNOR_1_1_NAND2_NUM200_OUT), .A2 (XNOR_1_2_NAND2_NUM200_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM200 (.ZN (N690), .A1 (XNOR_1_3_NAND2_NUM200_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM201_OUT, XNOR_1_2_NAND2_NUM201_OUT, XNOR_1_3_NAND2_NUM201_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM201 (.ZN (XNOR_1_1_NAND2_NUM201_OUT), .A1 (N607), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM201 (.ZN (XNOR_1_2_NAND2_NUM201_OUT), .A1 (GND), .A2 (N666));
      NOR2_X1 XNOR_1_3_NAND2_NUM201 (.ZN (XNOR_1_3_NAND2_NUM201_OUT), .A1 (XNOR_1_1_NAND2_NUM201_OUT), .A2 (XNOR_1_2_NAND2_NUM201_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM201 (.ZN (N691), .A1 (XNOR_1_3_NAND2_NUM201_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM202_OUT, XNOR_1_2_NAND2_NUM202_OUT, XNOR_1_3_NAND2_NUM202_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM202 (.ZN (XNOR_1_1_NAND2_NUM202_OUT), .A1 (N612), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM202 (.ZN (XNOR_1_2_NAND2_NUM202_OUT), .A1 (GND), .A2 (N669));
      NOR2_X1 XNOR_1_3_NAND2_NUM202 (.ZN (XNOR_1_3_NAND2_NUM202_OUT), .A1 (XNOR_1_1_NAND2_NUM202_OUT), .A2 (XNOR_1_2_NAND2_NUM202_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM202 (.ZN (N692), .A1 (XNOR_1_3_NAND2_NUM202_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM203_OUT, XNOR_1_2_NAND2_NUM203_OUT, XNOR_1_3_NAND2_NUM203_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM203 (.ZN (XNOR_1_1_NAND2_NUM203_OUT), .A1 (N617), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM203 (.ZN (XNOR_1_2_NAND2_NUM203_OUT), .A1 (GND), .A2 (N669));
      NOR2_X1 XNOR_1_3_NAND2_NUM203 (.ZN (XNOR_1_3_NAND2_NUM203_OUT), .A1 (XNOR_1_1_NAND2_NUM203_OUT), .A2 (XNOR_1_2_NAND2_NUM203_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM203 (.ZN (N693), .A1 (XNOR_1_3_NAND2_NUM203_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM204_OUT, XNOR_1_2_NAND2_NUM204_OUT, XNOR_1_3_NAND2_NUM204_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM204 (.ZN (XNOR_1_1_NAND2_NUM204_OUT), .A1 (N602), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM204 (.ZN (XNOR_1_2_NAND2_NUM204_OUT), .A1 (GND), .A2 (N672));
      NOR2_X1 XNOR_1_3_NAND2_NUM204 (.ZN (XNOR_1_3_NAND2_NUM204_OUT), .A1 (XNOR_1_1_NAND2_NUM204_OUT), .A2 (XNOR_1_2_NAND2_NUM204_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM204 (.ZN (N694), .A1 (XNOR_1_3_NAND2_NUM204_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM205_OUT, XNOR_1_2_NAND2_NUM205_OUT, XNOR_1_3_NAND2_NUM205_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM205 (.ZN (XNOR_1_1_NAND2_NUM205_OUT), .A1 (N612), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM205 (.ZN (XNOR_1_2_NAND2_NUM205_OUT), .A1 (GND), .A2 (N672));
      NOR2_X1 XNOR_1_3_NAND2_NUM205 (.ZN (XNOR_1_3_NAND2_NUM205_OUT), .A1 (XNOR_1_1_NAND2_NUM205_OUT), .A2 (XNOR_1_2_NAND2_NUM205_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM205 (.ZN (N695), .A1 (XNOR_1_3_NAND2_NUM205_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM206_OUT, XNOR_1_2_NAND2_NUM206_OUT, XNOR_1_3_NAND2_NUM206_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM206 (.ZN (XNOR_1_1_NAND2_NUM206_OUT), .A1 (N607), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM206 (.ZN (XNOR_1_2_NAND2_NUM206_OUT), .A1 (GND), .A2 (N675));
      NOR2_X1 XNOR_1_3_NAND2_NUM206 (.ZN (XNOR_1_3_NAND2_NUM206_OUT), .A1 (XNOR_1_1_NAND2_NUM206_OUT), .A2 (XNOR_1_2_NAND2_NUM206_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM206 (.ZN (N696), .A1 (XNOR_1_3_NAND2_NUM206_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM207_OUT, XNOR_1_2_NAND2_NUM207_OUT, XNOR_1_3_NAND2_NUM207_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM207 (.ZN (XNOR_1_1_NAND2_NUM207_OUT), .A1 (N617), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM207 (.ZN (XNOR_1_2_NAND2_NUM207_OUT), .A1 (GND), .A2 (N675));
      NOR2_X1 XNOR_1_3_NAND2_NUM207 (.ZN (XNOR_1_3_NAND2_NUM207_OUT), .A1 (XNOR_1_1_NAND2_NUM207_OUT), .A2 (XNOR_1_2_NAND2_NUM207_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM207 (.ZN (N697), .A1 (XNOR_1_3_NAND2_NUM207_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM208_OUT, XNOR_1_2_NAND2_NUM208_OUT, XNOR_1_3_NAND2_NUM208_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM208 (.ZN (XNOR_1_1_NAND2_NUM208_OUT), .A1 (N622), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM208 (.ZN (XNOR_1_2_NAND2_NUM208_OUT), .A1 (GND), .A2 (N678));
      NOR2_X1 XNOR_1_3_NAND2_NUM208 (.ZN (XNOR_1_3_NAND2_NUM208_OUT), .A1 (XNOR_1_1_NAND2_NUM208_OUT), .A2 (XNOR_1_2_NAND2_NUM208_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM208 (.ZN (N698), .A1 (XNOR_1_3_NAND2_NUM208_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM209_OUT, XNOR_1_2_NAND2_NUM209_OUT, XNOR_1_3_NAND2_NUM209_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM209 (.ZN (XNOR_1_1_NAND2_NUM209_OUT), .A1 (N627), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM209 (.ZN (XNOR_1_2_NAND2_NUM209_OUT), .A1 (GND), .A2 (N678));
      NOR2_X1 XNOR_1_3_NAND2_NUM209 (.ZN (XNOR_1_3_NAND2_NUM209_OUT), .A1 (XNOR_1_1_NAND2_NUM209_OUT), .A2 (XNOR_1_2_NAND2_NUM209_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM209 (.ZN (N699), .A1 (XNOR_1_3_NAND2_NUM209_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM210_OUT, XNOR_1_2_NAND2_NUM210_OUT, XNOR_1_3_NAND2_NUM210_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM210 (.ZN (XNOR_1_1_NAND2_NUM210_OUT), .A1 (N632), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM210 (.ZN (XNOR_1_2_NAND2_NUM210_OUT), .A1 (GND), .A2 (N681));
      NOR2_X1 XNOR_1_3_NAND2_NUM210 (.ZN (XNOR_1_3_NAND2_NUM210_OUT), .A1 (XNOR_1_1_NAND2_NUM210_OUT), .A2 (XNOR_1_2_NAND2_NUM210_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM210 (.ZN (N700), .A1 (XNOR_1_3_NAND2_NUM210_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM211_OUT, XNOR_1_2_NAND2_NUM211_OUT, XNOR_1_3_NAND2_NUM211_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM211 (.ZN (XNOR_1_1_NAND2_NUM211_OUT), .A1 (N637), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM211 (.ZN (XNOR_1_2_NAND2_NUM211_OUT), .A1 (GND), .A2 (N681));
      NOR2_X1 XNOR_1_3_NAND2_NUM211 (.ZN (XNOR_1_3_NAND2_NUM211_OUT), .A1 (XNOR_1_1_NAND2_NUM211_OUT), .A2 (XNOR_1_2_NAND2_NUM211_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM211 (.ZN (N701), .A1 (XNOR_1_3_NAND2_NUM211_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM212_OUT, XNOR_1_2_NAND2_NUM212_OUT, XNOR_1_3_NAND2_NUM212_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM212 (.ZN (XNOR_1_1_NAND2_NUM212_OUT), .A1 (N622), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM212 (.ZN (XNOR_1_2_NAND2_NUM212_OUT), .A1 (GND), .A2 (N684));
      NOR2_X1 XNOR_1_3_NAND2_NUM212 (.ZN (XNOR_1_3_NAND2_NUM212_OUT), .A1 (XNOR_1_1_NAND2_NUM212_OUT), .A2 (XNOR_1_2_NAND2_NUM212_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM212 (.ZN (N702), .A1 (XNOR_1_3_NAND2_NUM212_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM213_OUT, XNOR_1_2_NAND2_NUM213_OUT, XNOR_1_3_NAND2_NUM213_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM213 (.ZN (XNOR_1_1_NAND2_NUM213_OUT), .A1 (N632), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM213 (.ZN (XNOR_1_2_NAND2_NUM213_OUT), .A1 (GND), .A2 (N684));
      NOR2_X1 XNOR_1_3_NAND2_NUM213 (.ZN (XNOR_1_3_NAND2_NUM213_OUT), .A1 (XNOR_1_1_NAND2_NUM213_OUT), .A2 (XNOR_1_2_NAND2_NUM213_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM213 (.ZN (N703), .A1 (XNOR_1_3_NAND2_NUM213_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM214_OUT, XNOR_1_2_NAND2_NUM214_OUT, XNOR_1_3_NAND2_NUM214_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM214 (.ZN (XNOR_1_1_NAND2_NUM214_OUT), .A1 (N627), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM214 (.ZN (XNOR_1_2_NAND2_NUM214_OUT), .A1 (GND), .A2 (N687));
      NOR2_X1 XNOR_1_3_NAND2_NUM214 (.ZN (XNOR_1_3_NAND2_NUM214_OUT), .A1 (XNOR_1_1_NAND2_NUM214_OUT), .A2 (XNOR_1_2_NAND2_NUM214_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM214 (.ZN (N704), .A1 (XNOR_1_3_NAND2_NUM214_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM215_OUT, XNOR_1_2_NAND2_NUM215_OUT, XNOR_1_3_NAND2_NUM215_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM215 (.ZN (XNOR_1_1_NAND2_NUM215_OUT), .A1 (N637), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM215 (.ZN (XNOR_1_2_NAND2_NUM215_OUT), .A1 (GND), .A2 (N687));
      NOR2_X1 XNOR_1_3_NAND2_NUM215 (.ZN (XNOR_1_3_NAND2_NUM215_OUT), .A1 (XNOR_1_1_NAND2_NUM215_OUT), .A2 (XNOR_1_2_NAND2_NUM215_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM215 (.ZN (N705), .A1 (XNOR_1_3_NAND2_NUM215_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM216_OUT, XNOR_1_2_NAND2_NUM216_OUT, XNOR_1_3_NAND2_NUM216_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM216 (.ZN (XNOR_1_1_NAND2_NUM216_OUT), .A1 (N690), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM216 (.ZN (XNOR_1_2_NAND2_NUM216_OUT), .A1 (GND), .A2 (N691));
      NOR2_X1 XNOR_1_3_NAND2_NUM216 (.ZN (XNOR_1_3_NAND2_NUM216_OUT), .A1 (XNOR_1_1_NAND2_NUM216_OUT), .A2 (XNOR_1_2_NAND2_NUM216_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM216 (.ZN (N706), .A1 (XNOR_1_3_NAND2_NUM216_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM217_OUT, XNOR_1_2_NAND2_NUM217_OUT, XNOR_1_3_NAND2_NUM217_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM217 (.ZN (XNOR_1_1_NAND2_NUM217_OUT), .A1 (N692), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM217 (.ZN (XNOR_1_2_NAND2_NUM217_OUT), .A1 (GND), .A2 (N693));
      NOR2_X1 XNOR_1_3_NAND2_NUM217 (.ZN (XNOR_1_3_NAND2_NUM217_OUT), .A1 (XNOR_1_1_NAND2_NUM217_OUT), .A2 (XNOR_1_2_NAND2_NUM217_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM217 (.ZN (N709), .A1 (XNOR_1_3_NAND2_NUM217_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM218_OUT, XNOR_1_2_NAND2_NUM218_OUT, XNOR_1_3_NAND2_NUM218_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM218 (.ZN (XNOR_1_1_NAND2_NUM218_OUT), .A1 (N694), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM218 (.ZN (XNOR_1_2_NAND2_NUM218_OUT), .A1 (GND), .A2 (N695));
      NOR2_X1 XNOR_1_3_NAND2_NUM218 (.ZN (XNOR_1_3_NAND2_NUM218_OUT), .A1 (XNOR_1_1_NAND2_NUM218_OUT), .A2 (XNOR_1_2_NAND2_NUM218_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM218 (.ZN (N712), .A1 (XNOR_1_3_NAND2_NUM218_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM219_OUT, XNOR_1_2_NAND2_NUM219_OUT, XNOR_1_3_NAND2_NUM219_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM219 (.ZN (XNOR_1_1_NAND2_NUM219_OUT), .A1 (N696), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM219 (.ZN (XNOR_1_2_NAND2_NUM219_OUT), .A1 (GND), .A2 (N697));
      NOR2_X1 XNOR_1_3_NAND2_NUM219 (.ZN (XNOR_1_3_NAND2_NUM219_OUT), .A1 (XNOR_1_1_NAND2_NUM219_OUT), .A2 (XNOR_1_2_NAND2_NUM219_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM219 (.ZN (N715), .A1 (XNOR_1_3_NAND2_NUM219_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM220_OUT, XNOR_1_2_NAND2_NUM220_OUT, XNOR_1_3_NAND2_NUM220_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM220 (.ZN (XNOR_1_1_NAND2_NUM220_OUT), .A1 (N698), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM220 (.ZN (XNOR_1_2_NAND2_NUM220_OUT), .A1 (GND), .A2 (N699));
      NOR2_X1 XNOR_1_3_NAND2_NUM220 (.ZN (XNOR_1_3_NAND2_NUM220_OUT), .A1 (XNOR_1_1_NAND2_NUM220_OUT), .A2 (XNOR_1_2_NAND2_NUM220_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM220 (.ZN (N718), .A1 (XNOR_1_3_NAND2_NUM220_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM221_OUT, XNOR_1_2_NAND2_NUM221_OUT, XNOR_1_3_NAND2_NUM221_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM221 (.ZN (XNOR_1_1_NAND2_NUM221_OUT), .A1 (N700), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM221 (.ZN (XNOR_1_2_NAND2_NUM221_OUT), .A1 (GND), .A2 (N701));
      NOR2_X1 XNOR_1_3_NAND2_NUM221 (.ZN (XNOR_1_3_NAND2_NUM221_OUT), .A1 (XNOR_1_1_NAND2_NUM221_OUT), .A2 (XNOR_1_2_NAND2_NUM221_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM221 (.ZN (N721), .A1 (XNOR_1_3_NAND2_NUM221_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM222_OUT, XNOR_1_2_NAND2_NUM222_OUT, XNOR_1_3_NAND2_NUM222_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM222 (.ZN (XNOR_1_1_NAND2_NUM222_OUT), .A1 (N702), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM222 (.ZN (XNOR_1_2_NAND2_NUM222_OUT), .A1 (GND), .A2 (N703));
      NOR2_X1 XNOR_1_3_NAND2_NUM222 (.ZN (XNOR_1_3_NAND2_NUM222_OUT), .A1 (XNOR_1_1_NAND2_NUM222_OUT), .A2 (XNOR_1_2_NAND2_NUM222_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM222 (.ZN (N724), .A1 (XNOR_1_3_NAND2_NUM222_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM223_OUT, XNOR_1_2_NAND2_NUM223_OUT, XNOR_1_3_NAND2_NUM223_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM223 (.ZN (XNOR_1_1_NAND2_NUM223_OUT), .A1 (N704), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM223 (.ZN (XNOR_1_2_NAND2_NUM223_OUT), .A1 (GND), .A2 (N705));
      NOR2_X1 XNOR_1_3_NAND2_NUM223 (.ZN (XNOR_1_3_NAND2_NUM223_OUT), .A1 (XNOR_1_1_NAND2_NUM223_OUT), .A2 (XNOR_1_2_NAND2_NUM223_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM223 (.ZN (N727), .A1 (XNOR_1_3_NAND2_NUM223_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM224_OUT, XNOR_1_2_NAND2_NUM224_OUT, XNOR_1_3_NAND2_NUM224_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM224 (.ZN (XNOR_1_1_NAND2_NUM224_OUT), .A1 (N242), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM224 (.ZN (XNOR_1_2_NAND2_NUM224_OUT), .A1 (GND), .A2 (N718));
      NOR2_X1 XNOR_1_3_NAND2_NUM224 (.ZN (XNOR_1_3_NAND2_NUM224_OUT), .A1 (XNOR_1_1_NAND2_NUM224_OUT), .A2 (XNOR_1_2_NAND2_NUM224_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM224 (.ZN (N730), .A1 (XNOR_1_3_NAND2_NUM224_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM225_OUT, XNOR_1_2_NAND2_NUM225_OUT, XNOR_1_3_NAND2_NUM225_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM225 (.ZN (XNOR_1_1_NAND2_NUM225_OUT), .A1 (N245), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM225 (.ZN (XNOR_1_2_NAND2_NUM225_OUT), .A1 (GND), .A2 (N721));
      NOR2_X1 XNOR_1_3_NAND2_NUM225 (.ZN (XNOR_1_3_NAND2_NUM225_OUT), .A1 (XNOR_1_1_NAND2_NUM225_OUT), .A2 (XNOR_1_2_NAND2_NUM225_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM225 (.ZN (N733), .A1 (XNOR_1_3_NAND2_NUM225_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM226_OUT, XNOR_1_2_NAND2_NUM226_OUT, XNOR_1_3_NAND2_NUM226_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM226 (.ZN (XNOR_1_1_NAND2_NUM226_OUT), .A1 (N248), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM226 (.ZN (XNOR_1_2_NAND2_NUM226_OUT), .A1 (GND), .A2 (N724));
      NOR2_X1 XNOR_1_3_NAND2_NUM226 (.ZN (XNOR_1_3_NAND2_NUM226_OUT), .A1 (XNOR_1_1_NAND2_NUM226_OUT), .A2 (XNOR_1_2_NAND2_NUM226_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM226 (.ZN (N736), .A1 (XNOR_1_3_NAND2_NUM226_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM227_OUT, XNOR_1_2_NAND2_NUM227_OUT, XNOR_1_3_NAND2_NUM227_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM227 (.ZN (XNOR_1_1_NAND2_NUM227_OUT), .A1 (N251), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM227 (.ZN (XNOR_1_2_NAND2_NUM227_OUT), .A1 (GND), .A2 (N727));
      NOR2_X1 XNOR_1_3_NAND2_NUM227 (.ZN (XNOR_1_3_NAND2_NUM227_OUT), .A1 (XNOR_1_1_NAND2_NUM227_OUT), .A2 (XNOR_1_2_NAND2_NUM227_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM227 (.ZN (N739), .A1 (XNOR_1_3_NAND2_NUM227_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM228_OUT, XNOR_1_2_NAND2_NUM228_OUT, XNOR_1_3_NAND2_NUM228_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM228 (.ZN (XNOR_1_1_NAND2_NUM228_OUT), .A1 (N254), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM228 (.ZN (XNOR_1_2_NAND2_NUM228_OUT), .A1 (GND), .A2 (N706));
      NOR2_X1 XNOR_1_3_NAND2_NUM228 (.ZN (XNOR_1_3_NAND2_NUM228_OUT), .A1 (XNOR_1_1_NAND2_NUM228_OUT), .A2 (XNOR_1_2_NAND2_NUM228_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM228 (.ZN (N742), .A1 (XNOR_1_3_NAND2_NUM228_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM229_OUT, XNOR_1_2_NAND2_NUM229_OUT, XNOR_1_3_NAND2_NUM229_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM229 (.ZN (XNOR_1_1_NAND2_NUM229_OUT), .A1 (N257), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM229 (.ZN (XNOR_1_2_NAND2_NUM229_OUT), .A1 (GND), .A2 (N709));
      NOR2_X1 XNOR_1_3_NAND2_NUM229 (.ZN (XNOR_1_3_NAND2_NUM229_OUT), .A1 (XNOR_1_1_NAND2_NUM229_OUT), .A2 (XNOR_1_2_NAND2_NUM229_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM229 (.ZN (N745), .A1 (XNOR_1_3_NAND2_NUM229_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM230_OUT, XNOR_1_2_NAND2_NUM230_OUT, XNOR_1_3_NAND2_NUM230_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM230 (.ZN (XNOR_1_1_NAND2_NUM230_OUT), .A1 (N260), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM230 (.ZN (XNOR_1_2_NAND2_NUM230_OUT), .A1 (GND), .A2 (N712));
      NOR2_X1 XNOR_1_3_NAND2_NUM230 (.ZN (XNOR_1_3_NAND2_NUM230_OUT), .A1 (XNOR_1_1_NAND2_NUM230_OUT), .A2 (XNOR_1_2_NAND2_NUM230_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM230 (.ZN (N748), .A1 (XNOR_1_3_NAND2_NUM230_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM231_OUT, XNOR_1_2_NAND2_NUM231_OUT, XNOR_1_3_NAND2_NUM231_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM231 (.ZN (XNOR_1_1_NAND2_NUM231_OUT), .A1 (N263), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM231 (.ZN (XNOR_1_2_NAND2_NUM231_OUT), .A1 (GND), .A2 (N715));
      NOR2_X1 XNOR_1_3_NAND2_NUM231 (.ZN (XNOR_1_3_NAND2_NUM231_OUT), .A1 (XNOR_1_1_NAND2_NUM231_OUT), .A2 (XNOR_1_2_NAND2_NUM231_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM231 (.ZN (N751), .A1 (XNOR_1_3_NAND2_NUM231_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM232_OUT, XNOR_1_2_NAND2_NUM232_OUT, XNOR_1_3_NAND2_NUM232_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM232 (.ZN (XNOR_1_1_NAND2_NUM232_OUT), .A1 (N242), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM232 (.ZN (XNOR_1_2_NAND2_NUM232_OUT), .A1 (GND), .A2 (N730));
      NOR2_X1 XNOR_1_3_NAND2_NUM232 (.ZN (XNOR_1_3_NAND2_NUM232_OUT), .A1 (XNOR_1_1_NAND2_NUM232_OUT), .A2 (XNOR_1_2_NAND2_NUM232_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM232 (.ZN (N754), .A1 (XNOR_1_3_NAND2_NUM232_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM233_OUT, XNOR_1_2_NAND2_NUM233_OUT, XNOR_1_3_NAND2_NUM233_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM233 (.ZN (XNOR_1_1_NAND2_NUM233_OUT), .A1 (N718), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM233 (.ZN (XNOR_1_2_NAND2_NUM233_OUT), .A1 (GND), .A2 (N730));
      NOR2_X1 XNOR_1_3_NAND2_NUM233 (.ZN (XNOR_1_3_NAND2_NUM233_OUT), .A1 (XNOR_1_1_NAND2_NUM233_OUT), .A2 (XNOR_1_2_NAND2_NUM233_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM233 (.ZN (N755), .A1 (XNOR_1_3_NAND2_NUM233_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM234_OUT, XNOR_1_2_NAND2_NUM234_OUT, XNOR_1_3_NAND2_NUM234_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM234 (.ZN (XNOR_1_1_NAND2_NUM234_OUT), .A1 (N245), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM234 (.ZN (XNOR_1_2_NAND2_NUM234_OUT), .A1 (GND), .A2 (N733));
      NOR2_X1 XNOR_1_3_NAND2_NUM234 (.ZN (XNOR_1_3_NAND2_NUM234_OUT), .A1 (XNOR_1_1_NAND2_NUM234_OUT), .A2 (XNOR_1_2_NAND2_NUM234_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM234 (.ZN (N756), .A1 (XNOR_1_3_NAND2_NUM234_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM235_OUT, XNOR_1_2_NAND2_NUM235_OUT, XNOR_1_3_NAND2_NUM235_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM235 (.ZN (XNOR_1_1_NAND2_NUM235_OUT), .A1 (N721), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM235 (.ZN (XNOR_1_2_NAND2_NUM235_OUT), .A1 (GND), .A2 (N733));
      NOR2_X1 XNOR_1_3_NAND2_NUM235 (.ZN (XNOR_1_3_NAND2_NUM235_OUT), .A1 (XNOR_1_1_NAND2_NUM235_OUT), .A2 (XNOR_1_2_NAND2_NUM235_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM235 (.ZN (N757), .A1 (XNOR_1_3_NAND2_NUM235_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM236_OUT, XNOR_1_2_NAND2_NUM236_OUT, XNOR_1_3_NAND2_NUM236_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM236 (.ZN (XNOR_1_1_NAND2_NUM236_OUT), .A1 (N248), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM236 (.ZN (XNOR_1_2_NAND2_NUM236_OUT), .A1 (GND), .A2 (N736));
      NOR2_X1 XNOR_1_3_NAND2_NUM236 (.ZN (XNOR_1_3_NAND2_NUM236_OUT), .A1 (XNOR_1_1_NAND2_NUM236_OUT), .A2 (XNOR_1_2_NAND2_NUM236_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM236 (.ZN (N758), .A1 (XNOR_1_3_NAND2_NUM236_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM237_OUT, XNOR_1_2_NAND2_NUM237_OUT, XNOR_1_3_NAND2_NUM237_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM237 (.ZN (XNOR_1_1_NAND2_NUM237_OUT), .A1 (N724), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM237 (.ZN (XNOR_1_2_NAND2_NUM237_OUT), .A1 (GND), .A2 (N736));
      NOR2_X1 XNOR_1_3_NAND2_NUM237 (.ZN (XNOR_1_3_NAND2_NUM237_OUT), .A1 (XNOR_1_1_NAND2_NUM237_OUT), .A2 (XNOR_1_2_NAND2_NUM237_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM237 (.ZN (N759), .A1 (XNOR_1_3_NAND2_NUM237_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM238_OUT, XNOR_1_2_NAND2_NUM238_OUT, XNOR_1_3_NAND2_NUM238_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM238 (.ZN (XNOR_1_1_NAND2_NUM238_OUT), .A1 (N251), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM238 (.ZN (XNOR_1_2_NAND2_NUM238_OUT), .A1 (GND), .A2 (N739));
      NOR2_X1 XNOR_1_3_NAND2_NUM238 (.ZN (XNOR_1_3_NAND2_NUM238_OUT), .A1 (XNOR_1_1_NAND2_NUM238_OUT), .A2 (XNOR_1_2_NAND2_NUM238_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM238 (.ZN (N760), .A1 (XNOR_1_3_NAND2_NUM238_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM239_OUT, XNOR_1_2_NAND2_NUM239_OUT, XNOR_1_3_NAND2_NUM239_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM239 (.ZN (XNOR_1_1_NAND2_NUM239_OUT), .A1 (N727), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM239 (.ZN (XNOR_1_2_NAND2_NUM239_OUT), .A1 (GND), .A2 (N739));
      NOR2_X1 XNOR_1_3_NAND2_NUM239 (.ZN (XNOR_1_3_NAND2_NUM239_OUT), .A1 (XNOR_1_1_NAND2_NUM239_OUT), .A2 (XNOR_1_2_NAND2_NUM239_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM239 (.ZN (N761), .A1 (XNOR_1_3_NAND2_NUM239_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM240_OUT, XNOR_1_2_NAND2_NUM240_OUT, XNOR_1_3_NAND2_NUM240_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM240 (.ZN (XNOR_1_1_NAND2_NUM240_OUT), .A1 (N254), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM240 (.ZN (XNOR_1_2_NAND2_NUM240_OUT), .A1 (GND), .A2 (N742));
      NOR2_X1 XNOR_1_3_NAND2_NUM240 (.ZN (XNOR_1_3_NAND2_NUM240_OUT), .A1 (XNOR_1_1_NAND2_NUM240_OUT), .A2 (XNOR_1_2_NAND2_NUM240_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM240 (.ZN (N762), .A1 (XNOR_1_3_NAND2_NUM240_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM241_OUT, XNOR_1_2_NAND2_NUM241_OUT, XNOR_1_3_NAND2_NUM241_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM241 (.ZN (XNOR_1_1_NAND2_NUM241_OUT), .A1 (N706), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM241 (.ZN (XNOR_1_2_NAND2_NUM241_OUT), .A1 (GND), .A2 (N742));
      NOR2_X1 XNOR_1_3_NAND2_NUM241 (.ZN (XNOR_1_3_NAND2_NUM241_OUT), .A1 (XNOR_1_1_NAND2_NUM241_OUT), .A2 (XNOR_1_2_NAND2_NUM241_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM241 (.ZN (N763), .A1 (XNOR_1_3_NAND2_NUM241_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM242_OUT, XNOR_1_2_NAND2_NUM242_OUT, XNOR_1_3_NAND2_NUM242_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM242 (.ZN (XNOR_1_1_NAND2_NUM242_OUT), .A1 (N257), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM242 (.ZN (XNOR_1_2_NAND2_NUM242_OUT), .A1 (GND), .A2 (N745));
      NOR2_X1 XNOR_1_3_NAND2_NUM242 (.ZN (XNOR_1_3_NAND2_NUM242_OUT), .A1 (XNOR_1_1_NAND2_NUM242_OUT), .A2 (XNOR_1_2_NAND2_NUM242_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM242 (.ZN (N764), .A1 (XNOR_1_3_NAND2_NUM242_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM243_OUT, XNOR_1_2_NAND2_NUM243_OUT, XNOR_1_3_NAND2_NUM243_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM243 (.ZN (XNOR_1_1_NAND2_NUM243_OUT), .A1 (N709), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM243 (.ZN (XNOR_1_2_NAND2_NUM243_OUT), .A1 (GND), .A2 (N745));
      NOR2_X1 XNOR_1_3_NAND2_NUM243 (.ZN (XNOR_1_3_NAND2_NUM243_OUT), .A1 (XNOR_1_1_NAND2_NUM243_OUT), .A2 (XNOR_1_2_NAND2_NUM243_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM243 (.ZN (N765), .A1 (XNOR_1_3_NAND2_NUM243_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM244_OUT, XNOR_1_2_NAND2_NUM244_OUT, XNOR_1_3_NAND2_NUM244_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM244 (.ZN (XNOR_1_1_NAND2_NUM244_OUT), .A1 (N260), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM244 (.ZN (XNOR_1_2_NAND2_NUM244_OUT), .A1 (GND), .A2 (N748));
      NOR2_X1 XNOR_1_3_NAND2_NUM244 (.ZN (XNOR_1_3_NAND2_NUM244_OUT), .A1 (XNOR_1_1_NAND2_NUM244_OUT), .A2 (XNOR_1_2_NAND2_NUM244_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM244 (.ZN (N766), .A1 (XNOR_1_3_NAND2_NUM244_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM245_OUT, XNOR_1_2_NAND2_NUM245_OUT, XNOR_1_3_NAND2_NUM245_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM245 (.ZN (XNOR_1_1_NAND2_NUM245_OUT), .A1 (N712), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM245 (.ZN (XNOR_1_2_NAND2_NUM245_OUT), .A1 (GND), .A2 (N748));
      NOR2_X1 XNOR_1_3_NAND2_NUM245 (.ZN (XNOR_1_3_NAND2_NUM245_OUT), .A1 (XNOR_1_1_NAND2_NUM245_OUT), .A2 (XNOR_1_2_NAND2_NUM245_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM245 (.ZN (N767), .A1 (XNOR_1_3_NAND2_NUM245_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM246_OUT, XNOR_1_2_NAND2_NUM246_OUT, XNOR_1_3_NAND2_NUM246_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM246 (.ZN (XNOR_1_1_NAND2_NUM246_OUT), .A1 (N263), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM246 (.ZN (XNOR_1_2_NAND2_NUM246_OUT), .A1 (GND), .A2 (N751));
      NOR2_X1 XNOR_1_3_NAND2_NUM246 (.ZN (XNOR_1_3_NAND2_NUM246_OUT), .A1 (XNOR_1_1_NAND2_NUM246_OUT), .A2 (XNOR_1_2_NAND2_NUM246_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM246 (.ZN (N768), .A1 (XNOR_1_3_NAND2_NUM246_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM247_OUT, XNOR_1_2_NAND2_NUM247_OUT, XNOR_1_3_NAND2_NUM247_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM247 (.ZN (XNOR_1_1_NAND2_NUM247_OUT), .A1 (N715), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM247 (.ZN (XNOR_1_2_NAND2_NUM247_OUT), .A1 (GND), .A2 (N751));
      NOR2_X1 XNOR_1_3_NAND2_NUM247 (.ZN (XNOR_1_3_NAND2_NUM247_OUT), .A1 (XNOR_1_1_NAND2_NUM247_OUT), .A2 (XNOR_1_2_NAND2_NUM247_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM247 (.ZN (N769), .A1 (XNOR_1_3_NAND2_NUM247_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM248_OUT, XNOR_1_2_NAND2_NUM248_OUT, XNOR_1_3_NAND2_NUM248_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM248 (.ZN (XNOR_1_1_NAND2_NUM248_OUT), .A1 (N754), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM248 (.ZN (XNOR_1_2_NAND2_NUM248_OUT), .A1 (GND), .A2 (N755));
      NOR2_X1 XNOR_1_3_NAND2_NUM248 (.ZN (XNOR_1_3_NAND2_NUM248_OUT), .A1 (XNOR_1_1_NAND2_NUM248_OUT), .A2 (XNOR_1_2_NAND2_NUM248_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM248 (.ZN (N770), .A1 (XNOR_1_3_NAND2_NUM248_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM249_OUT, XNOR_1_2_NAND2_NUM249_OUT, XNOR_1_3_NAND2_NUM249_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM249 (.ZN (XNOR_1_1_NAND2_NUM249_OUT), .A1 (N756), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM249 (.ZN (XNOR_1_2_NAND2_NUM249_OUT), .A1 (GND), .A2 (N757));
      NOR2_X1 XNOR_1_3_NAND2_NUM249 (.ZN (XNOR_1_3_NAND2_NUM249_OUT), .A1 (XNOR_1_1_NAND2_NUM249_OUT), .A2 (XNOR_1_2_NAND2_NUM249_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM249 (.ZN (N773), .A1 (XNOR_1_3_NAND2_NUM249_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM250_OUT, XNOR_1_2_NAND2_NUM250_OUT, XNOR_1_3_NAND2_NUM250_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM250 (.ZN (XNOR_1_1_NAND2_NUM250_OUT), .A1 (N758), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM250 (.ZN (XNOR_1_2_NAND2_NUM250_OUT), .A1 (GND), .A2 (N759));
      NOR2_X1 XNOR_1_3_NAND2_NUM250 (.ZN (XNOR_1_3_NAND2_NUM250_OUT), .A1 (XNOR_1_1_NAND2_NUM250_OUT), .A2 (XNOR_1_2_NAND2_NUM250_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM250 (.ZN (N776), .A1 (XNOR_1_3_NAND2_NUM250_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM251_OUT, XNOR_1_2_NAND2_NUM251_OUT, XNOR_1_3_NAND2_NUM251_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM251 (.ZN (XNOR_1_1_NAND2_NUM251_OUT), .A1 (N760), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM251 (.ZN (XNOR_1_2_NAND2_NUM251_OUT), .A1 (GND), .A2 (N761));
      NOR2_X1 XNOR_1_3_NAND2_NUM251 (.ZN (XNOR_1_3_NAND2_NUM251_OUT), .A1 (XNOR_1_1_NAND2_NUM251_OUT), .A2 (XNOR_1_2_NAND2_NUM251_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM251 (.ZN (N779), .A1 (XNOR_1_3_NAND2_NUM251_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM252_OUT, XNOR_1_2_NAND2_NUM252_OUT, XNOR_1_3_NAND2_NUM252_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM252 (.ZN (XNOR_1_1_NAND2_NUM252_OUT), .A1 (N762), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM252 (.ZN (XNOR_1_2_NAND2_NUM252_OUT), .A1 (GND), .A2 (N763));
      NOR2_X1 XNOR_1_3_NAND2_NUM252 (.ZN (XNOR_1_3_NAND2_NUM252_OUT), .A1 (XNOR_1_1_NAND2_NUM252_OUT), .A2 (XNOR_1_2_NAND2_NUM252_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM252 (.ZN (N782), .A1 (XNOR_1_3_NAND2_NUM252_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM253_OUT, XNOR_1_2_NAND2_NUM253_OUT, XNOR_1_3_NAND2_NUM253_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM253 (.ZN (XNOR_1_1_NAND2_NUM253_OUT), .A1 (N764), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM253 (.ZN (XNOR_1_2_NAND2_NUM253_OUT), .A1 (GND), .A2 (N765));
      NOR2_X1 XNOR_1_3_NAND2_NUM253 (.ZN (XNOR_1_3_NAND2_NUM253_OUT), .A1 (XNOR_1_1_NAND2_NUM253_OUT), .A2 (XNOR_1_2_NAND2_NUM253_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM253 (.ZN (N785), .A1 (XNOR_1_3_NAND2_NUM253_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM254_OUT, XNOR_1_2_NAND2_NUM254_OUT, XNOR_1_3_NAND2_NUM254_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM254 (.ZN (XNOR_1_1_NAND2_NUM254_OUT), .A1 (N766), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM254 (.ZN (XNOR_1_2_NAND2_NUM254_OUT), .A1 (GND), .A2 (N767));
      NOR2_X1 XNOR_1_3_NAND2_NUM254 (.ZN (XNOR_1_3_NAND2_NUM254_OUT), .A1 (XNOR_1_1_NAND2_NUM254_OUT), .A2 (XNOR_1_2_NAND2_NUM254_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM254 (.ZN (N788), .A1 (XNOR_1_3_NAND2_NUM254_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM255_OUT, XNOR_1_2_NAND2_NUM255_OUT, XNOR_1_3_NAND2_NUM255_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM255 (.ZN (XNOR_1_1_NAND2_NUM255_OUT), .A1 (N768), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM255 (.ZN (XNOR_1_2_NAND2_NUM255_OUT), .A1 (GND), .A2 (N769));
      NOR2_X1 XNOR_1_3_NAND2_NUM255 (.ZN (XNOR_1_3_NAND2_NUM255_OUT), .A1 (XNOR_1_1_NAND2_NUM255_OUT), .A2 (XNOR_1_2_NAND2_NUM255_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM255 (.ZN (N791), .A1 (XNOR_1_3_NAND2_NUM255_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM256_OUT, XNOR_1_2_NAND2_NUM256_OUT, XNOR_1_3_NAND2_NUM256_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM256 (.ZN (XNOR_1_1_NAND2_NUM256_OUT), .A1 (N642), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM256 (.ZN (XNOR_1_2_NAND2_NUM256_OUT), .A1 (GND), .A2 (N770));
      NOR2_X1 XNOR_1_3_NAND2_NUM256 (.ZN (XNOR_1_3_NAND2_NUM256_OUT), .A1 (XNOR_1_1_NAND2_NUM256_OUT), .A2 (XNOR_1_2_NAND2_NUM256_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM256 (.ZN (N794), .A1 (XNOR_1_3_NAND2_NUM256_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM257_OUT, XNOR_1_2_NAND2_NUM257_OUT, XNOR_1_3_NAND2_NUM257_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM257 (.ZN (XNOR_1_1_NAND2_NUM257_OUT), .A1 (N645), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM257 (.ZN (XNOR_1_2_NAND2_NUM257_OUT), .A1 (GND), .A2 (N773));
      NOR2_X1 XNOR_1_3_NAND2_NUM257 (.ZN (XNOR_1_3_NAND2_NUM257_OUT), .A1 (XNOR_1_1_NAND2_NUM257_OUT), .A2 (XNOR_1_2_NAND2_NUM257_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM257 (.ZN (N797), .A1 (XNOR_1_3_NAND2_NUM257_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM258_OUT, XNOR_1_2_NAND2_NUM258_OUT, XNOR_1_3_NAND2_NUM258_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM258 (.ZN (XNOR_1_1_NAND2_NUM258_OUT), .A1 (N648), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM258 (.ZN (XNOR_1_2_NAND2_NUM258_OUT), .A1 (GND), .A2 (N776));
      NOR2_X1 XNOR_1_3_NAND2_NUM258 (.ZN (XNOR_1_3_NAND2_NUM258_OUT), .A1 (XNOR_1_1_NAND2_NUM258_OUT), .A2 (XNOR_1_2_NAND2_NUM258_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM258 (.ZN (N800), .A1 (XNOR_1_3_NAND2_NUM258_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM259_OUT, XNOR_1_2_NAND2_NUM259_OUT, XNOR_1_3_NAND2_NUM259_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM259 (.ZN (XNOR_1_1_NAND2_NUM259_OUT), .A1 (N651), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM259 (.ZN (XNOR_1_2_NAND2_NUM259_OUT), .A1 (GND), .A2 (N779));
      NOR2_X1 XNOR_1_3_NAND2_NUM259 (.ZN (XNOR_1_3_NAND2_NUM259_OUT), .A1 (XNOR_1_1_NAND2_NUM259_OUT), .A2 (XNOR_1_2_NAND2_NUM259_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM259 (.ZN (N803), .A1 (XNOR_1_3_NAND2_NUM259_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM260_OUT, XNOR_1_2_NAND2_NUM260_OUT, XNOR_1_3_NAND2_NUM260_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM260 (.ZN (XNOR_1_1_NAND2_NUM260_OUT), .A1 (N654), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM260 (.ZN (XNOR_1_2_NAND2_NUM260_OUT), .A1 (GND), .A2 (N782));
      NOR2_X1 XNOR_1_3_NAND2_NUM260 (.ZN (XNOR_1_3_NAND2_NUM260_OUT), .A1 (XNOR_1_1_NAND2_NUM260_OUT), .A2 (XNOR_1_2_NAND2_NUM260_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM260 (.ZN (N806), .A1 (XNOR_1_3_NAND2_NUM260_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM261_OUT, XNOR_1_2_NAND2_NUM261_OUT, XNOR_1_3_NAND2_NUM261_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM261 (.ZN (XNOR_1_1_NAND2_NUM261_OUT), .A1 (N657), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM261 (.ZN (XNOR_1_2_NAND2_NUM261_OUT), .A1 (GND), .A2 (N785));
      NOR2_X1 XNOR_1_3_NAND2_NUM261 (.ZN (XNOR_1_3_NAND2_NUM261_OUT), .A1 (XNOR_1_1_NAND2_NUM261_OUT), .A2 (XNOR_1_2_NAND2_NUM261_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM261 (.ZN (N809), .A1 (XNOR_1_3_NAND2_NUM261_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM262_OUT, XNOR_1_2_NAND2_NUM262_OUT, XNOR_1_3_NAND2_NUM262_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM262 (.ZN (XNOR_1_1_NAND2_NUM262_OUT), .A1 (N660), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM262 (.ZN (XNOR_1_2_NAND2_NUM262_OUT), .A1 (GND), .A2 (N788));
      NOR2_X1 XNOR_1_3_NAND2_NUM262 (.ZN (XNOR_1_3_NAND2_NUM262_OUT), .A1 (XNOR_1_1_NAND2_NUM262_OUT), .A2 (XNOR_1_2_NAND2_NUM262_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM262 (.ZN (N812), .A1 (XNOR_1_3_NAND2_NUM262_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM263_OUT, XNOR_1_2_NAND2_NUM263_OUT, XNOR_1_3_NAND2_NUM263_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM263 (.ZN (XNOR_1_1_NAND2_NUM263_OUT), .A1 (N663), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM263 (.ZN (XNOR_1_2_NAND2_NUM263_OUT), .A1 (GND), .A2 (N791));
      NOR2_X1 XNOR_1_3_NAND2_NUM263 (.ZN (XNOR_1_3_NAND2_NUM263_OUT), .A1 (XNOR_1_1_NAND2_NUM263_OUT), .A2 (XNOR_1_2_NAND2_NUM263_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM263 (.ZN (N815), .A1 (XNOR_1_3_NAND2_NUM263_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM264_OUT, XNOR_1_2_NAND2_NUM264_OUT, XNOR_1_3_NAND2_NUM264_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM264 (.ZN (XNOR_1_1_NAND2_NUM264_OUT), .A1 (N642), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM264 (.ZN (XNOR_1_2_NAND2_NUM264_OUT), .A1 (GND), .A2 (N794));
      NOR2_X1 XNOR_1_3_NAND2_NUM264 (.ZN (XNOR_1_3_NAND2_NUM264_OUT), .A1 (XNOR_1_1_NAND2_NUM264_OUT), .A2 (XNOR_1_2_NAND2_NUM264_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM264 (.ZN (N818), .A1 (XNOR_1_3_NAND2_NUM264_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM265_OUT, XNOR_1_2_NAND2_NUM265_OUT, XNOR_1_3_NAND2_NUM265_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM265 (.ZN (XNOR_1_1_NAND2_NUM265_OUT), .A1 (N770), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM265 (.ZN (XNOR_1_2_NAND2_NUM265_OUT), .A1 (GND), .A2 (N794));
      NOR2_X1 XNOR_1_3_NAND2_NUM265 (.ZN (XNOR_1_3_NAND2_NUM265_OUT), .A1 (XNOR_1_1_NAND2_NUM265_OUT), .A2 (XNOR_1_2_NAND2_NUM265_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM265 (.ZN (N819), .A1 (XNOR_1_3_NAND2_NUM265_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM266_OUT, XNOR_1_2_NAND2_NUM266_OUT, XNOR_1_3_NAND2_NUM266_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM266 (.ZN (XNOR_1_1_NAND2_NUM266_OUT), .A1 (N645), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM266 (.ZN (XNOR_1_2_NAND2_NUM266_OUT), .A1 (GND), .A2 (N797));
      NOR2_X1 XNOR_1_3_NAND2_NUM266 (.ZN (XNOR_1_3_NAND2_NUM266_OUT), .A1 (XNOR_1_1_NAND2_NUM266_OUT), .A2 (XNOR_1_2_NAND2_NUM266_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM266 (.ZN (N820), .A1 (XNOR_1_3_NAND2_NUM266_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM267_OUT, XNOR_1_2_NAND2_NUM267_OUT, XNOR_1_3_NAND2_NUM267_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM267 (.ZN (XNOR_1_1_NAND2_NUM267_OUT), .A1 (N773), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM267 (.ZN (XNOR_1_2_NAND2_NUM267_OUT), .A1 (GND), .A2 (N797));
      NOR2_X1 XNOR_1_3_NAND2_NUM267 (.ZN (XNOR_1_3_NAND2_NUM267_OUT), .A1 (XNOR_1_1_NAND2_NUM267_OUT), .A2 (XNOR_1_2_NAND2_NUM267_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM267 (.ZN (N821), .A1 (XNOR_1_3_NAND2_NUM267_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM268_OUT, XNOR_1_2_NAND2_NUM268_OUT, XNOR_1_3_NAND2_NUM268_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM268 (.ZN (XNOR_1_1_NAND2_NUM268_OUT), .A1 (N648), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM268 (.ZN (XNOR_1_2_NAND2_NUM268_OUT), .A1 (GND), .A2 (N800));
      NOR2_X1 XNOR_1_3_NAND2_NUM268 (.ZN (XNOR_1_3_NAND2_NUM268_OUT), .A1 (XNOR_1_1_NAND2_NUM268_OUT), .A2 (XNOR_1_2_NAND2_NUM268_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM268 (.ZN (N822), .A1 (XNOR_1_3_NAND2_NUM268_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM269_OUT, XNOR_1_2_NAND2_NUM269_OUT, XNOR_1_3_NAND2_NUM269_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM269 (.ZN (XNOR_1_1_NAND2_NUM269_OUT), .A1 (N776), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM269 (.ZN (XNOR_1_2_NAND2_NUM269_OUT), .A1 (GND), .A2 (N800));
      NOR2_X1 XNOR_1_3_NAND2_NUM269 (.ZN (XNOR_1_3_NAND2_NUM269_OUT), .A1 (XNOR_1_1_NAND2_NUM269_OUT), .A2 (XNOR_1_2_NAND2_NUM269_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM269 (.ZN (N823), .A1 (XNOR_1_3_NAND2_NUM269_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM270_OUT, XNOR_1_2_NAND2_NUM270_OUT, XNOR_1_3_NAND2_NUM270_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM270 (.ZN (XNOR_1_1_NAND2_NUM270_OUT), .A1 (N651), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM270 (.ZN (XNOR_1_2_NAND2_NUM270_OUT), .A1 (GND), .A2 (N803));
      NOR2_X1 XNOR_1_3_NAND2_NUM270 (.ZN (XNOR_1_3_NAND2_NUM270_OUT), .A1 (XNOR_1_1_NAND2_NUM270_OUT), .A2 (XNOR_1_2_NAND2_NUM270_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM270 (.ZN (N824), .A1 (XNOR_1_3_NAND2_NUM270_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM271_OUT, XNOR_1_2_NAND2_NUM271_OUT, XNOR_1_3_NAND2_NUM271_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM271 (.ZN (XNOR_1_1_NAND2_NUM271_OUT), .A1 (N779), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM271 (.ZN (XNOR_1_2_NAND2_NUM271_OUT), .A1 (GND), .A2 (N803));
      NOR2_X1 XNOR_1_3_NAND2_NUM271 (.ZN (XNOR_1_3_NAND2_NUM271_OUT), .A1 (XNOR_1_1_NAND2_NUM271_OUT), .A2 (XNOR_1_2_NAND2_NUM271_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM271 (.ZN (N825), .A1 (XNOR_1_3_NAND2_NUM271_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM272_OUT, XNOR_1_2_NAND2_NUM272_OUT, XNOR_1_3_NAND2_NUM272_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM272 (.ZN (XNOR_1_1_NAND2_NUM272_OUT), .A1 (N654), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM272 (.ZN (XNOR_1_2_NAND2_NUM272_OUT), .A1 (GND), .A2 (N806));
      NOR2_X1 XNOR_1_3_NAND2_NUM272 (.ZN (XNOR_1_3_NAND2_NUM272_OUT), .A1 (XNOR_1_1_NAND2_NUM272_OUT), .A2 (XNOR_1_2_NAND2_NUM272_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM272 (.ZN (N826), .A1 (XNOR_1_3_NAND2_NUM272_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM273_OUT, XNOR_1_2_NAND2_NUM273_OUT, XNOR_1_3_NAND2_NUM273_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM273 (.ZN (XNOR_1_1_NAND2_NUM273_OUT), .A1 (N782), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM273 (.ZN (XNOR_1_2_NAND2_NUM273_OUT), .A1 (GND), .A2 (N806));
      NOR2_X1 XNOR_1_3_NAND2_NUM273 (.ZN (XNOR_1_3_NAND2_NUM273_OUT), .A1 (XNOR_1_1_NAND2_NUM273_OUT), .A2 (XNOR_1_2_NAND2_NUM273_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM273 (.ZN (N827), .A1 (XNOR_1_3_NAND2_NUM273_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM274_OUT, XNOR_1_2_NAND2_NUM274_OUT, XNOR_1_3_NAND2_NUM274_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM274 (.ZN (XNOR_1_1_NAND2_NUM274_OUT), .A1 (N657), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM274 (.ZN (XNOR_1_2_NAND2_NUM274_OUT), .A1 (GND), .A2 (N809));
      NOR2_X1 XNOR_1_3_NAND2_NUM274 (.ZN (XNOR_1_3_NAND2_NUM274_OUT), .A1 (XNOR_1_1_NAND2_NUM274_OUT), .A2 (XNOR_1_2_NAND2_NUM274_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM274 (.ZN (N828), .A1 (XNOR_1_3_NAND2_NUM274_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM275_OUT, XNOR_1_2_NAND2_NUM275_OUT, XNOR_1_3_NAND2_NUM275_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM275 (.ZN (XNOR_1_1_NAND2_NUM275_OUT), .A1 (N785), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM275 (.ZN (XNOR_1_2_NAND2_NUM275_OUT), .A1 (GND), .A2 (N809));
      NOR2_X1 XNOR_1_3_NAND2_NUM275 (.ZN (XNOR_1_3_NAND2_NUM275_OUT), .A1 (XNOR_1_1_NAND2_NUM275_OUT), .A2 (XNOR_1_2_NAND2_NUM275_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM275 (.ZN (N829), .A1 (XNOR_1_3_NAND2_NUM275_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM276_OUT, XNOR_1_2_NAND2_NUM276_OUT, XNOR_1_3_NAND2_NUM276_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM276 (.ZN (XNOR_1_1_NAND2_NUM276_OUT), .A1 (N660), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM276 (.ZN (XNOR_1_2_NAND2_NUM276_OUT), .A1 (GND), .A2 (N812));
      NOR2_X1 XNOR_1_3_NAND2_NUM276 (.ZN (XNOR_1_3_NAND2_NUM276_OUT), .A1 (XNOR_1_1_NAND2_NUM276_OUT), .A2 (XNOR_1_2_NAND2_NUM276_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM276 (.ZN (N830), .A1 (XNOR_1_3_NAND2_NUM276_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM277_OUT, XNOR_1_2_NAND2_NUM277_OUT, XNOR_1_3_NAND2_NUM277_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM277 (.ZN (XNOR_1_1_NAND2_NUM277_OUT), .A1 (N788), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM277 (.ZN (XNOR_1_2_NAND2_NUM277_OUT), .A1 (GND), .A2 (N812));
      NOR2_X1 XNOR_1_3_NAND2_NUM277 (.ZN (XNOR_1_3_NAND2_NUM277_OUT), .A1 (XNOR_1_1_NAND2_NUM277_OUT), .A2 (XNOR_1_2_NAND2_NUM277_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM277 (.ZN (N831), .A1 (XNOR_1_3_NAND2_NUM277_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM278_OUT, XNOR_1_2_NAND2_NUM278_OUT, XNOR_1_3_NAND2_NUM278_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM278 (.ZN (XNOR_1_1_NAND2_NUM278_OUT), .A1 (N663), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM278 (.ZN (XNOR_1_2_NAND2_NUM278_OUT), .A1 (GND), .A2 (N815));
      NOR2_X1 XNOR_1_3_NAND2_NUM278 (.ZN (XNOR_1_3_NAND2_NUM278_OUT), .A1 (XNOR_1_1_NAND2_NUM278_OUT), .A2 (XNOR_1_2_NAND2_NUM278_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM278 (.ZN (N832), .A1 (XNOR_1_3_NAND2_NUM278_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM279_OUT, XNOR_1_2_NAND2_NUM279_OUT, XNOR_1_3_NAND2_NUM279_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM279 (.ZN (XNOR_1_1_NAND2_NUM279_OUT), .A1 (N791), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM279 (.ZN (XNOR_1_2_NAND2_NUM279_OUT), .A1 (GND), .A2 (N815));
      NOR2_X1 XNOR_1_3_NAND2_NUM279 (.ZN (XNOR_1_3_NAND2_NUM279_OUT), .A1 (XNOR_1_1_NAND2_NUM279_OUT), .A2 (XNOR_1_2_NAND2_NUM279_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM279 (.ZN (N833), .A1 (XNOR_1_3_NAND2_NUM279_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM280_OUT, XNOR_1_2_NAND2_NUM280_OUT, XNOR_1_3_NAND2_NUM280_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM280 (.ZN (XNOR_1_1_NAND2_NUM280_OUT), .A1 (N818), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM280 (.ZN (XNOR_1_2_NAND2_NUM280_OUT), .A1 (GND), .A2 (N819));
      NOR2_X1 XNOR_1_3_NAND2_NUM280 (.ZN (XNOR_1_3_NAND2_NUM280_OUT), .A1 (XNOR_1_1_NAND2_NUM280_OUT), .A2 (XNOR_1_2_NAND2_NUM280_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM280 (.ZN (N834), .A1 (XNOR_1_3_NAND2_NUM280_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM281_OUT, XNOR_1_2_NAND2_NUM281_OUT, XNOR_1_3_NAND2_NUM281_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM281 (.ZN (XNOR_1_1_NAND2_NUM281_OUT), .A1 (N820), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM281 (.ZN (XNOR_1_2_NAND2_NUM281_OUT), .A1 (GND), .A2 (N821));
      NOR2_X1 XNOR_1_3_NAND2_NUM281 (.ZN (XNOR_1_3_NAND2_NUM281_OUT), .A1 (XNOR_1_1_NAND2_NUM281_OUT), .A2 (XNOR_1_2_NAND2_NUM281_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM281 (.ZN (N847), .A1 (XNOR_1_3_NAND2_NUM281_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM282_OUT, XNOR_1_2_NAND2_NUM282_OUT, XNOR_1_3_NAND2_NUM282_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM282 (.ZN (XNOR_1_1_NAND2_NUM282_OUT), .A1 (N822), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM282 (.ZN (XNOR_1_2_NAND2_NUM282_OUT), .A1 (GND), .A2 (N823));
      NOR2_X1 XNOR_1_3_NAND2_NUM282 (.ZN (XNOR_1_3_NAND2_NUM282_OUT), .A1 (XNOR_1_1_NAND2_NUM282_OUT), .A2 (XNOR_1_2_NAND2_NUM282_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM282 (.ZN (N860), .A1 (XNOR_1_3_NAND2_NUM282_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM283_OUT, XNOR_1_2_NAND2_NUM283_OUT, XNOR_1_3_NAND2_NUM283_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM283 (.ZN (XNOR_1_1_NAND2_NUM283_OUT), .A1 (N824), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM283 (.ZN (XNOR_1_2_NAND2_NUM283_OUT), .A1 (GND), .A2 (N825));
      NOR2_X1 XNOR_1_3_NAND2_NUM283 (.ZN (XNOR_1_3_NAND2_NUM283_OUT), .A1 (XNOR_1_1_NAND2_NUM283_OUT), .A2 (XNOR_1_2_NAND2_NUM283_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM283 (.ZN (N873), .A1 (XNOR_1_3_NAND2_NUM283_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM284_OUT, XNOR_1_2_NAND2_NUM284_OUT, XNOR_1_3_NAND2_NUM284_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM284 (.ZN (XNOR_1_1_NAND2_NUM284_OUT), .A1 (N828), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM284 (.ZN (XNOR_1_2_NAND2_NUM284_OUT), .A1 (GND), .A2 (N829));
      NOR2_X1 XNOR_1_3_NAND2_NUM284 (.ZN (XNOR_1_3_NAND2_NUM284_OUT), .A1 (XNOR_1_1_NAND2_NUM284_OUT), .A2 (XNOR_1_2_NAND2_NUM284_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM284 (.ZN (N886), .A1 (XNOR_1_3_NAND2_NUM284_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM285_OUT, XNOR_1_2_NAND2_NUM285_OUT, XNOR_1_3_NAND2_NUM285_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM285 (.ZN (XNOR_1_1_NAND2_NUM285_OUT), .A1 (N832), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM285 (.ZN (XNOR_1_2_NAND2_NUM285_OUT), .A1 (GND), .A2 (N833));
      NOR2_X1 XNOR_1_3_NAND2_NUM285 (.ZN (XNOR_1_3_NAND2_NUM285_OUT), .A1 (XNOR_1_1_NAND2_NUM285_OUT), .A2 (XNOR_1_2_NAND2_NUM285_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM285 (.ZN (N899), .A1 (XNOR_1_3_NAND2_NUM285_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM286_OUT, XNOR_1_2_NAND2_NUM286_OUT, XNOR_1_3_NAND2_NUM286_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM286 (.ZN (XNOR_1_1_NAND2_NUM286_OUT), .A1 (N830), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM286 (.ZN (XNOR_1_2_NAND2_NUM286_OUT), .A1 (GND), .A2 (N831));
      NOR2_X1 XNOR_1_3_NAND2_NUM286 (.ZN (XNOR_1_3_NAND2_NUM286_OUT), .A1 (XNOR_1_1_NAND2_NUM286_OUT), .A2 (XNOR_1_2_NAND2_NUM286_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM286 (.ZN (N912), .A1 (XNOR_1_3_NAND2_NUM286_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM287_OUT, XNOR_1_2_NAND2_NUM287_OUT, XNOR_1_3_NAND2_NUM287_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM287 (.ZN (XNOR_1_1_NAND2_NUM287_OUT), .A1 (N826), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM287 (.ZN (XNOR_1_2_NAND2_NUM287_OUT), .A1 (GND), .A2 (N827));
      NOR2_X1 XNOR_1_3_NAND2_NUM287 (.ZN (XNOR_1_3_NAND2_NUM287_OUT), .A1 (XNOR_1_1_NAND2_NUM287_OUT), .A2 (XNOR_1_2_NAND2_NUM287_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM287 (.ZN (N925), .A1 (XNOR_1_3_NAND2_NUM287_OUT), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM0 (.ZN (N938), .A1 (N834), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM1 (.ZN (N939), .A1 (N847), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM2 (.ZN (N940), .A1 (N860), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM3 (.ZN (N941), .A1 (N834), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM4 (.ZN (N942), .A1 (N847), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM5 (.ZN (N943), .A1 (N873), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM6 (.ZN (N944), .A1 (N834), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM7 (.ZN (N945), .A1 (N860), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM8 (.ZN (N946), .A1 (N873), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM9 (.ZN (N947), .A1 (N847), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM10 (.ZN (N948), .A1 (N860), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM11 (.ZN (N949), .A1 (N873), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM12 (.ZN (N950), .A1 (N886), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM13 (.ZN (N951), .A1 (N899), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM14 (.ZN (N952), .A1 (N886), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM15 (.ZN (N953), .A1 (N912), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM16 (.ZN (N954), .A1 (N925), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM17 (.ZN (N955), .A1 (N899), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM18 (.ZN (N956), .A1 (N925), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM19 (.ZN (N957), .A1 (N912), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM20 (.ZN (N958), .A1 (N925), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM21 (.ZN (N959), .A1 (N886), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM22 (.ZN (N960), .A1 (N912), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM23 (.ZN (N961), .A1 (N925), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM24 (.ZN (N962), .A1 (N886), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM25 (.ZN (N963), .A1 (N899), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM26 (.ZN (N964), .A1 (N925), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM27 (.ZN (N965), .A1 (N912), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM28 (.ZN (N966), .A1 (N899), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM29 (.ZN (N967), .A1 (N886), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM30 (.ZN (N968), .A1 (N912), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM31 (.ZN (N969), .A1 (N899), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM32 (.ZN (N970), .A1 (N847), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM33 (.ZN (N971), .A1 (N873), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM34 (.ZN (N972), .A1 (N847), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM35 (.ZN (N973), .A1 (N860), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM36 (.ZN (N974), .A1 (N834), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM37 (.ZN (N975), .A1 (N873), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM38 (.ZN (N976), .A1 (N834), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM39 (.ZN (N977), .A1 (N860), .A2 (GND));
      wire XNOR_1_1_AND4_NUM0_OUT, XNOR_1_2_AND4_NUM0_OUT, XNOR_1_3_AND4_NUM0_OUT;
      NOR2_X1 XNOR_1_1_AND4_NUM0 (.ZN (XNOR_1_1_AND4_NUM0_OUT), .A1 (N938), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND4_NUM0 (.ZN (XNOR_1_2_AND4_NUM0_OUT), .A1 (GND), .A2 (N939));
      NOR2_X1 XNOR_1_3_AND4_NUM0 (.ZN (XNOR_1_3_AND4_NUM0_OUT), .A1 (XNOR_1_1_AND4_NUM0_OUT), .A2 (XNOR_1_2_AND4_NUM0_OUT));

      wire XNOR_2_1_AND4_NUM0_OUT, XNOR_2_2_AND4_NUM0_OUT, XNOR_2_3_AND4_NUM0_OUT;
      NOR2_X1 XNOR_2_1_AND4_NUM0 (.ZN (XNOR_2_1_AND4_NUM0_OUT), .A1 (N940), .A2 (GND));
      NOR2_X1 XNOR_2_2_AND4_NUM0 (.ZN (XNOR_2_2_AND4_NUM0_OUT), .A1 (GND), .A2 (N873));
      NOR2_X1 XNOR_2_3_AND4_NUM0 (.ZN (XNOR_2_3_AND4_NUM0_OUT), .A1 (XNOR_2_1_AND4_NUM0_OUT), .A2 (XNOR_2_2_AND4_NUM0_OUT));

      wire XNOR_3_1_AND4_NUM0_OUT, XNOR_3_2_AND4_NUM0_OUT;
      NOR2_X1 XNOR_3_1_AND4_NUM0 (.ZN (XNOR_3_1_AND4_NUM0_OUT), .A1 (XNOR_1_3_AND4_NUM0_OUT), .A2 (GND));
      NOR2_X1 XNOR_3_2_AND4_NUM0 (.ZN (XNOR_3_2_AND4_NUM0_OUT), .A1 (GND), .A2 (XNOR_2_3_AND4_NUM0_OUT));
      NOR2_X1 XNOR_3_3_AND4_NUM0 (.ZN (N978), .A1 (XNOR_3_1_AND4_NUM0_OUT), .A2 (XNOR_3_2_AND4_NUM0_OUT));
      wire XNOR_1_1_AND4_NUM1_OUT, XNOR_1_2_AND4_NUM1_OUT, XNOR_1_3_AND4_NUM1_OUT;
      NOR2_X1 XNOR_1_1_AND4_NUM1 (.ZN (XNOR_1_1_AND4_NUM1_OUT), .A1 (N941), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND4_NUM1 (.ZN (XNOR_1_2_AND4_NUM1_OUT), .A1 (GND), .A2 (N942));
      NOR2_X1 XNOR_1_3_AND4_NUM1 (.ZN (XNOR_1_3_AND4_NUM1_OUT), .A1 (XNOR_1_1_AND4_NUM1_OUT), .A2 (XNOR_1_2_AND4_NUM1_OUT));

      wire XNOR_2_1_AND4_NUM1_OUT, XNOR_2_2_AND4_NUM1_OUT, XNOR_2_3_AND4_NUM1_OUT;
      NOR2_X1 XNOR_2_1_AND4_NUM1 (.ZN (XNOR_2_1_AND4_NUM1_OUT), .A1 (N860), .A2 (GND));
      NOR2_X1 XNOR_2_2_AND4_NUM1 (.ZN (XNOR_2_2_AND4_NUM1_OUT), .A1 (GND), .A2 (N943));
      NOR2_X1 XNOR_2_3_AND4_NUM1 (.ZN (XNOR_2_3_AND4_NUM1_OUT), .A1 (XNOR_2_1_AND4_NUM1_OUT), .A2 (XNOR_2_2_AND4_NUM1_OUT));

      wire XNOR_3_1_AND4_NUM1_OUT, XNOR_3_2_AND4_NUM1_OUT;
      NOR2_X1 XNOR_3_1_AND4_NUM1 (.ZN (XNOR_3_1_AND4_NUM1_OUT), .A1 (XNOR_1_3_AND4_NUM1_OUT), .A2 (GND));
      NOR2_X1 XNOR_3_2_AND4_NUM1 (.ZN (XNOR_3_2_AND4_NUM1_OUT), .A1 (GND), .A2 (XNOR_2_3_AND4_NUM1_OUT));
      NOR2_X1 XNOR_3_3_AND4_NUM1 (.ZN (N979), .A1 (XNOR_3_1_AND4_NUM1_OUT), .A2 (XNOR_3_2_AND4_NUM1_OUT));
      wire XNOR_1_1_AND4_NUM2_OUT, XNOR_1_2_AND4_NUM2_OUT, XNOR_1_3_AND4_NUM2_OUT;
      NOR2_X1 XNOR_1_1_AND4_NUM2 (.ZN (XNOR_1_1_AND4_NUM2_OUT), .A1 (N944), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND4_NUM2 (.ZN (XNOR_1_2_AND4_NUM2_OUT), .A1 (GND), .A2 (N847));
      NOR2_X1 XNOR_1_3_AND4_NUM2 (.ZN (XNOR_1_3_AND4_NUM2_OUT), .A1 (XNOR_1_1_AND4_NUM2_OUT), .A2 (XNOR_1_2_AND4_NUM2_OUT));

      wire XNOR_2_1_AND4_NUM2_OUT, XNOR_2_2_AND4_NUM2_OUT, XNOR_2_3_AND4_NUM2_OUT;
      NOR2_X1 XNOR_2_1_AND4_NUM2 (.ZN (XNOR_2_1_AND4_NUM2_OUT), .A1 (N945), .A2 (GND));
      NOR2_X1 XNOR_2_2_AND4_NUM2 (.ZN (XNOR_2_2_AND4_NUM2_OUT), .A1 (GND), .A2 (N946));
      NOR2_X1 XNOR_2_3_AND4_NUM2 (.ZN (XNOR_2_3_AND4_NUM2_OUT), .A1 (XNOR_2_1_AND4_NUM2_OUT), .A2 (XNOR_2_2_AND4_NUM2_OUT));

      wire XNOR_3_1_AND4_NUM2_OUT, XNOR_3_2_AND4_NUM2_OUT;
      NOR2_X1 XNOR_3_1_AND4_NUM2 (.ZN (XNOR_3_1_AND4_NUM2_OUT), .A1 (XNOR_1_3_AND4_NUM2_OUT), .A2 (GND));
      NOR2_X1 XNOR_3_2_AND4_NUM2 (.ZN (XNOR_3_2_AND4_NUM2_OUT), .A1 (GND), .A2 (XNOR_2_3_AND4_NUM2_OUT));
      NOR2_X1 XNOR_3_3_AND4_NUM2 (.ZN (N980), .A1 (XNOR_3_1_AND4_NUM2_OUT), .A2 (XNOR_3_2_AND4_NUM2_OUT));
      wire XNOR_1_1_AND4_NUM3_OUT, XNOR_1_2_AND4_NUM3_OUT, XNOR_1_3_AND4_NUM3_OUT;
      NOR2_X1 XNOR_1_1_AND4_NUM3 (.ZN (XNOR_1_1_AND4_NUM3_OUT), .A1 (N834), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND4_NUM3 (.ZN (XNOR_1_2_AND4_NUM3_OUT), .A1 (GND), .A2 (N947));
      NOR2_X1 XNOR_1_3_AND4_NUM3 (.ZN (XNOR_1_3_AND4_NUM3_OUT), .A1 (XNOR_1_1_AND4_NUM3_OUT), .A2 (XNOR_1_2_AND4_NUM3_OUT));

      wire XNOR_2_1_AND4_NUM3_OUT, XNOR_2_2_AND4_NUM3_OUT, XNOR_2_3_AND4_NUM3_OUT;
      NOR2_X1 XNOR_2_1_AND4_NUM3 (.ZN (XNOR_2_1_AND4_NUM3_OUT), .A1 (N948), .A2 (GND));
      NOR2_X1 XNOR_2_2_AND4_NUM3 (.ZN (XNOR_2_2_AND4_NUM3_OUT), .A1 (GND), .A2 (N949));
      NOR2_X1 XNOR_2_3_AND4_NUM3 (.ZN (XNOR_2_3_AND4_NUM3_OUT), .A1 (XNOR_2_1_AND4_NUM3_OUT), .A2 (XNOR_2_2_AND4_NUM3_OUT));

      wire XNOR_3_1_AND4_NUM3_OUT, XNOR_3_2_AND4_NUM3_OUT;
      NOR2_X1 XNOR_3_1_AND4_NUM3 (.ZN (XNOR_3_1_AND4_NUM3_OUT), .A1 (XNOR_1_3_AND4_NUM3_OUT), .A2 (GND));
      NOR2_X1 XNOR_3_2_AND4_NUM3 (.ZN (XNOR_3_2_AND4_NUM3_OUT), .A1 (GND), .A2 (XNOR_2_3_AND4_NUM3_OUT));
      NOR2_X1 XNOR_3_3_AND4_NUM3 (.ZN (N981), .A1 (XNOR_3_1_AND4_NUM3_OUT), .A2 (XNOR_3_2_AND4_NUM3_OUT));
      wire XNOR_1_1_AND4_NUM4_OUT, XNOR_1_2_AND4_NUM4_OUT, XNOR_1_3_AND4_NUM4_OUT;
      NOR2_X1 XNOR_1_1_AND4_NUM4 (.ZN (XNOR_1_1_AND4_NUM4_OUT), .A1 (N958), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND4_NUM4 (.ZN (XNOR_1_2_AND4_NUM4_OUT), .A1 (GND), .A2 (N959));
      NOR2_X1 XNOR_1_3_AND4_NUM4 (.ZN (XNOR_1_3_AND4_NUM4_OUT), .A1 (XNOR_1_1_AND4_NUM4_OUT), .A2 (XNOR_1_2_AND4_NUM4_OUT));

      wire XNOR_2_1_AND4_NUM4_OUT, XNOR_2_2_AND4_NUM4_OUT, XNOR_2_3_AND4_NUM4_OUT;
      NOR2_X1 XNOR_2_1_AND4_NUM4 (.ZN (XNOR_2_1_AND4_NUM4_OUT), .A1 (N960), .A2 (GND));
      NOR2_X1 XNOR_2_2_AND4_NUM4 (.ZN (XNOR_2_2_AND4_NUM4_OUT), .A1 (GND), .A2 (N899));
      NOR2_X1 XNOR_2_3_AND4_NUM4 (.ZN (XNOR_2_3_AND4_NUM4_OUT), .A1 (XNOR_2_1_AND4_NUM4_OUT), .A2 (XNOR_2_2_AND4_NUM4_OUT));

      wire XNOR_3_1_AND4_NUM4_OUT, XNOR_3_2_AND4_NUM4_OUT;
      NOR2_X1 XNOR_3_1_AND4_NUM4 (.ZN (XNOR_3_1_AND4_NUM4_OUT), .A1 (XNOR_1_3_AND4_NUM4_OUT), .A2 (GND));
      NOR2_X1 XNOR_3_2_AND4_NUM4 (.ZN (XNOR_3_2_AND4_NUM4_OUT), .A1 (GND), .A2 (XNOR_2_3_AND4_NUM4_OUT));
      NOR2_X1 XNOR_3_3_AND4_NUM4 (.ZN (N982), .A1 (XNOR_3_1_AND4_NUM4_OUT), .A2 (XNOR_3_2_AND4_NUM4_OUT));
      wire XNOR_1_1_AND4_NUM5_OUT, XNOR_1_2_AND4_NUM5_OUT, XNOR_1_3_AND4_NUM5_OUT;
      NOR2_X1 XNOR_1_1_AND4_NUM5 (.ZN (XNOR_1_1_AND4_NUM5_OUT), .A1 (N961), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND4_NUM5 (.ZN (XNOR_1_2_AND4_NUM5_OUT), .A1 (GND), .A2 (N962));
      NOR2_X1 XNOR_1_3_AND4_NUM5 (.ZN (XNOR_1_3_AND4_NUM5_OUT), .A1 (XNOR_1_1_AND4_NUM5_OUT), .A2 (XNOR_1_2_AND4_NUM5_OUT));

      wire XNOR_2_1_AND4_NUM5_OUT, XNOR_2_2_AND4_NUM5_OUT, XNOR_2_3_AND4_NUM5_OUT;
      NOR2_X1 XNOR_2_1_AND4_NUM5 (.ZN (XNOR_2_1_AND4_NUM5_OUT), .A1 (N912), .A2 (GND));
      NOR2_X1 XNOR_2_2_AND4_NUM5 (.ZN (XNOR_2_2_AND4_NUM5_OUT), .A1 (GND), .A2 (N963));
      NOR2_X1 XNOR_2_3_AND4_NUM5 (.ZN (XNOR_2_3_AND4_NUM5_OUT), .A1 (XNOR_2_1_AND4_NUM5_OUT), .A2 (XNOR_2_2_AND4_NUM5_OUT));

      wire XNOR_3_1_AND4_NUM5_OUT, XNOR_3_2_AND4_NUM5_OUT;
      NOR2_X1 XNOR_3_1_AND4_NUM5 (.ZN (XNOR_3_1_AND4_NUM5_OUT), .A1 (XNOR_1_3_AND4_NUM5_OUT), .A2 (GND));
      NOR2_X1 XNOR_3_2_AND4_NUM5 (.ZN (XNOR_3_2_AND4_NUM5_OUT), .A1 (GND), .A2 (XNOR_2_3_AND4_NUM5_OUT));
      NOR2_X1 XNOR_3_3_AND4_NUM5 (.ZN (N983), .A1 (XNOR_3_1_AND4_NUM5_OUT), .A2 (XNOR_3_2_AND4_NUM5_OUT));
      wire XNOR_1_1_AND4_NUM6_OUT, XNOR_1_2_AND4_NUM6_OUT, XNOR_1_3_AND4_NUM6_OUT;
      NOR2_X1 XNOR_1_1_AND4_NUM6 (.ZN (XNOR_1_1_AND4_NUM6_OUT), .A1 (N964), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND4_NUM6 (.ZN (XNOR_1_2_AND4_NUM6_OUT), .A1 (GND), .A2 (N886));
      NOR2_X1 XNOR_1_3_AND4_NUM6 (.ZN (XNOR_1_3_AND4_NUM6_OUT), .A1 (XNOR_1_1_AND4_NUM6_OUT), .A2 (XNOR_1_2_AND4_NUM6_OUT));

      wire XNOR_2_1_AND4_NUM6_OUT, XNOR_2_2_AND4_NUM6_OUT, XNOR_2_3_AND4_NUM6_OUT;
      NOR2_X1 XNOR_2_1_AND4_NUM6 (.ZN (XNOR_2_1_AND4_NUM6_OUT), .A1 (N965), .A2 (GND));
      NOR2_X1 XNOR_2_2_AND4_NUM6 (.ZN (XNOR_2_2_AND4_NUM6_OUT), .A1 (GND), .A2 (N966));
      NOR2_X1 XNOR_2_3_AND4_NUM6 (.ZN (XNOR_2_3_AND4_NUM6_OUT), .A1 (XNOR_2_1_AND4_NUM6_OUT), .A2 (XNOR_2_2_AND4_NUM6_OUT));

      wire XNOR_3_1_AND4_NUM6_OUT, XNOR_3_2_AND4_NUM6_OUT;
      NOR2_X1 XNOR_3_1_AND4_NUM6 (.ZN (XNOR_3_1_AND4_NUM6_OUT), .A1 (XNOR_1_3_AND4_NUM6_OUT), .A2 (GND));
      NOR2_X1 XNOR_3_2_AND4_NUM6 (.ZN (XNOR_3_2_AND4_NUM6_OUT), .A1 (GND), .A2 (XNOR_2_3_AND4_NUM6_OUT));
      NOR2_X1 XNOR_3_3_AND4_NUM6 (.ZN (N984), .A1 (XNOR_3_1_AND4_NUM6_OUT), .A2 (XNOR_3_2_AND4_NUM6_OUT));
      wire XNOR_1_1_AND4_NUM7_OUT, XNOR_1_2_AND4_NUM7_OUT, XNOR_1_3_AND4_NUM7_OUT;
      NOR2_X1 XNOR_1_1_AND4_NUM7 (.ZN (XNOR_1_1_AND4_NUM7_OUT), .A1 (N925), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND4_NUM7 (.ZN (XNOR_1_2_AND4_NUM7_OUT), .A1 (GND), .A2 (N967));
      NOR2_X1 XNOR_1_3_AND4_NUM7 (.ZN (XNOR_1_3_AND4_NUM7_OUT), .A1 (XNOR_1_1_AND4_NUM7_OUT), .A2 (XNOR_1_2_AND4_NUM7_OUT));

      wire XNOR_2_1_AND4_NUM7_OUT, XNOR_2_2_AND4_NUM7_OUT, XNOR_2_3_AND4_NUM7_OUT;
      NOR2_X1 XNOR_2_1_AND4_NUM7 (.ZN (XNOR_2_1_AND4_NUM7_OUT), .A1 (N968), .A2 (GND));
      NOR2_X1 XNOR_2_2_AND4_NUM7 (.ZN (XNOR_2_2_AND4_NUM7_OUT), .A1 (GND), .A2 (N969));
      NOR2_X1 XNOR_2_3_AND4_NUM7 (.ZN (XNOR_2_3_AND4_NUM7_OUT), .A1 (XNOR_2_1_AND4_NUM7_OUT), .A2 (XNOR_2_2_AND4_NUM7_OUT));

      wire XNOR_3_1_AND4_NUM7_OUT, XNOR_3_2_AND4_NUM7_OUT;
      NOR2_X1 XNOR_3_1_AND4_NUM7 (.ZN (XNOR_3_1_AND4_NUM7_OUT), .A1 (XNOR_1_3_AND4_NUM7_OUT), .A2 (GND));
      NOR2_X1 XNOR_3_2_AND4_NUM7 (.ZN (XNOR_3_2_AND4_NUM7_OUT), .A1 (GND), .A2 (XNOR_2_3_AND4_NUM7_OUT));
      NOR2_X1 XNOR_3_3_AND4_NUM7 (.ZN (N985), .A1 (XNOR_3_1_AND4_NUM7_OUT), .A2 (XNOR_3_2_AND4_NUM7_OUT));
      wire XNOR_1_1_OR4_NUM0_OUT, XNOR_1_2_OR4_NUM0_OUT, XNOR_2_1_OR4_NUM0_OUT, XNOR_2_2_OR4_NUM0_OUT, XNOR_3_1_OR4_NUM0_OUT;
      NOR2_X1 XNOR_1_1_OR4_NUM0 (.ZN (XNOR_1_1_OR4_NUM0_OUT), .A1 (N978), .A2 (N979));
      NOR2_X1 XNOR_1_2_OR4_NUM0 (.ZN (XNOR_1_2_OR4_NUM0_OUT), .A1 (XNOR_1_1_OR4_NUM0_OUT), .A2 (GND));

      NOR2_X1 XNOR_2_1_OR4_NUM0 (.ZN (XNOR_2_1_OR4_NUM0_OUT), .A1 (N980), .A2 (N981));
      NOR2_X1 XNOR_2_2_OR4_NUM0 (.ZN (XNOR_2_2_OR4_NUM0_OUT), .A1 (XNOR_2_1_OR4_NUM0_OUT), .A2 (GND));

      NOR2_X1 XNOR_3_1_OR4_NUM0 (.ZN (XNOR_3_1_OR4_NUM0_OUT), .A1 (XNOR_1_2_OR4_NUM0_OUT), .A2 (XNOR_2_2_OR4_NUM0_OUT));
      NOR2_X1 XNOR_3_2_OR4_NUM0 (.ZN (N986), .A1 (XNOR_3_1_OR4_NUM0_OUT), .A2 (GND));
      wire XNOR_1_1_OR4_NUM1_OUT, XNOR_1_2_OR4_NUM1_OUT, XNOR_2_1_OR4_NUM1_OUT, XNOR_2_2_OR4_NUM1_OUT, XNOR_3_1_OR4_NUM1_OUT;
      NOR2_X1 XNOR_1_1_OR4_NUM1 (.ZN (XNOR_1_1_OR4_NUM1_OUT), .A1 (N982), .A2 (N983));
      NOR2_X1 XNOR_1_2_OR4_NUM1 (.ZN (XNOR_1_2_OR4_NUM1_OUT), .A1 (XNOR_1_1_OR4_NUM1_OUT), .A2 (GND));

      NOR2_X1 XNOR_2_1_OR4_NUM1 (.ZN (XNOR_2_1_OR4_NUM1_OUT), .A1 (N984), .A2 (N985));
      NOR2_X1 XNOR_2_2_OR4_NUM1 (.ZN (XNOR_2_2_OR4_NUM1_OUT), .A1 (XNOR_2_1_OR4_NUM1_OUT), .A2 (GND));

      NOR2_X1 XNOR_3_1_OR4_NUM1 (.ZN (XNOR_3_1_OR4_NUM1_OUT), .A1 (XNOR_1_2_OR4_NUM1_OUT), .A2 (XNOR_2_2_OR4_NUM1_OUT));
      NOR2_X1 XNOR_3_2_OR4_NUM1 (.ZN (N991), .A1 (XNOR_3_1_OR4_NUM1_OUT), .A2 (GND));
      wire XNOR_1_1_AND5_NUM0_OUT, XNOR_1_2_AND5_NUM0_OUT, XNOR_1_3_AND5_NUM0_OUT;
      NOR2_X1 XNOR_1_1_AND5_NUM0 (.ZN (XNOR_1_1_AND5_NUM0_OUT), .A1 (N925), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND5_NUM0 (.ZN (XNOR_1_2_AND5_NUM0_OUT), .A1 (GND), .A2 (N950));
      NOR2_X1 XNOR_1_3_AND5_NUM0 (.ZN (XNOR_1_3_AND5_NUM0_OUT), .A1 (XNOR_1_1_AND5_NUM0_OUT), .A2 (XNOR_1_2_AND5_NUM0_OUT));

      wire XNOR_2_1_AND5_NUM0_OUT, XNOR_2_2_AND5_NUM0_OUT, XNOR_2_3_AND5_NUM0_OUT;
      NOR2_X1 XNOR_2_1_AND5_NUM0 (.ZN (XNOR_2_1_AND5_NUM0_OUT), .A1 (N912), .A2 (GND));
      NOR2_X1 XNOR_2_2_AND5_NUM0 (.ZN (XNOR_2_2_AND5_NUM0_OUT), .A1 (GND), .A2 (N951));
      NOR2_X1 XNOR_2_3_AND5_NUM0 (.ZN (XNOR_2_3_AND5_NUM0_OUT), .A1 (XNOR_2_1_AND5_NUM0_OUT), .A2 (XNOR_2_2_AND5_NUM0_OUT));

      wire XNOR_3_1_AND5_NUM0_OUT, XNOR_3_2_AND5_NUM0_OUT, XNOR_3_3_AND5_NUM0_OUT;
      NOR2_X1 XNOR_3_1_AND5_NUM0 (.ZN (XNOR_3_1_AND5_NUM0_OUT), .A1 (XNOR_1_3_AND5_NUM0_OUT), .A2 (GND));
      NOR2_X1 XNOR_3_2_AND5_NUM0 (.ZN (XNOR_3_2_AND5_NUM0_OUT), .A1 (GND), .A2 (XNOR_2_3_AND5_NUM0_OUT));
      NOR2_X1 XNOR_3_3_AND5_NUM0 (.ZN (XNOR_3_3_AND5_NUM0_OUT), .A1 (XNOR_3_1_AND5_NUM0_OUT), .A2 (XNOR_3_2_AND5_NUM0_OUT));

      wire XNOR_4_1_AND5_NUM0_OUT, XNOR_4_2_AND5_NUM0_OUT;
      NOR2_X1 XNOR_4_1_AND5_NUM0 (.ZN (XNOR_4_1_AND5_NUM0_OUT), .A1 (N986), .A2 (GND));
      NOR2_X1 XNOR_4_2_AND5_NUM0 (.ZN (XNOR_4_2_AND5_NUM0_OUT), .A1 (GND), .A2 (XNOR_3_3_AND5_NUM0_OUT));
      NOR2_X1 XNOR_4_3_AND5_NUM0 (.ZN (N996), .A1 (XNOR_4_1_AND5_NUM0_OUT), .A2 (XNOR_4_2_AND5_NUM0_OUT));
      wire XNOR_1_1_AND5_NUM1_OUT, XNOR_1_2_AND5_NUM1_OUT, XNOR_1_3_AND5_NUM1_OUT;
      NOR2_X1 XNOR_1_1_AND5_NUM1 (.ZN (XNOR_1_1_AND5_NUM1_OUT), .A1 (N925), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND5_NUM1 (.ZN (XNOR_1_2_AND5_NUM1_OUT), .A1 (GND), .A2 (N952));
      NOR2_X1 XNOR_1_3_AND5_NUM1 (.ZN (XNOR_1_3_AND5_NUM1_OUT), .A1 (XNOR_1_1_AND5_NUM1_OUT), .A2 (XNOR_1_2_AND5_NUM1_OUT));

      wire XNOR_2_1_AND5_NUM1_OUT, XNOR_2_2_AND5_NUM1_OUT, XNOR_2_3_AND5_NUM1_OUT;
      NOR2_X1 XNOR_2_1_AND5_NUM1 (.ZN (XNOR_2_1_AND5_NUM1_OUT), .A1 (N953), .A2 (GND));
      NOR2_X1 XNOR_2_2_AND5_NUM1 (.ZN (XNOR_2_2_AND5_NUM1_OUT), .A1 (GND), .A2 (N899));
      NOR2_X1 XNOR_2_3_AND5_NUM1 (.ZN (XNOR_2_3_AND5_NUM1_OUT), .A1 (XNOR_2_1_AND5_NUM1_OUT), .A2 (XNOR_2_2_AND5_NUM1_OUT));

      wire XNOR_3_1_AND5_NUM1_OUT, XNOR_3_2_AND5_NUM1_OUT, XNOR_3_3_AND5_NUM1_OUT;
      NOR2_X1 XNOR_3_1_AND5_NUM1 (.ZN (XNOR_3_1_AND5_NUM1_OUT), .A1 (XNOR_1_3_AND5_NUM1_OUT), .A2 (GND));
      NOR2_X1 XNOR_3_2_AND5_NUM1 (.ZN (XNOR_3_2_AND5_NUM1_OUT), .A1 (GND), .A2 (XNOR_2_3_AND5_NUM1_OUT));
      NOR2_X1 XNOR_3_3_AND5_NUM1 (.ZN (XNOR_3_3_AND5_NUM1_OUT), .A1 (XNOR_3_1_AND5_NUM1_OUT), .A2 (XNOR_3_2_AND5_NUM1_OUT));

      wire XNOR_4_1_AND5_NUM1_OUT, XNOR_4_2_AND5_NUM1_OUT;
      NOR2_X1 XNOR_4_1_AND5_NUM1 (.ZN (XNOR_4_1_AND5_NUM1_OUT), .A1 (N986), .A2 (GND));
      NOR2_X1 XNOR_4_2_AND5_NUM1 (.ZN (XNOR_4_2_AND5_NUM1_OUT), .A1 (GND), .A2 (XNOR_3_3_AND5_NUM1_OUT));
      NOR2_X1 XNOR_4_3_AND5_NUM1 (.ZN (N1001), .A1 (XNOR_4_1_AND5_NUM1_OUT), .A2 (XNOR_4_2_AND5_NUM1_OUT));
      wire XNOR_1_1_AND5_NUM2_OUT, XNOR_1_2_AND5_NUM2_OUT, XNOR_1_3_AND5_NUM2_OUT;
      NOR2_X1 XNOR_1_1_AND5_NUM2 (.ZN (XNOR_1_1_AND5_NUM2_OUT), .A1 (N954), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND5_NUM2 (.ZN (XNOR_1_2_AND5_NUM2_OUT), .A1 (GND), .A2 (N886));
      NOR2_X1 XNOR_1_3_AND5_NUM2 (.ZN (XNOR_1_3_AND5_NUM2_OUT), .A1 (XNOR_1_1_AND5_NUM2_OUT), .A2 (XNOR_1_2_AND5_NUM2_OUT));

      wire XNOR_2_1_AND5_NUM2_OUT, XNOR_2_2_AND5_NUM2_OUT, XNOR_2_3_AND5_NUM2_OUT;
      NOR2_X1 XNOR_2_1_AND5_NUM2 (.ZN (XNOR_2_1_AND5_NUM2_OUT), .A1 (N912), .A2 (GND));
      NOR2_X1 XNOR_2_2_AND5_NUM2 (.ZN (XNOR_2_2_AND5_NUM2_OUT), .A1 (GND), .A2 (N955));
      NOR2_X1 XNOR_2_3_AND5_NUM2 (.ZN (XNOR_2_3_AND5_NUM2_OUT), .A1 (XNOR_2_1_AND5_NUM2_OUT), .A2 (XNOR_2_2_AND5_NUM2_OUT));

      wire XNOR_3_1_AND5_NUM2_OUT, XNOR_3_2_AND5_NUM2_OUT, XNOR_3_3_AND5_NUM2_OUT;
      NOR2_X1 XNOR_3_1_AND5_NUM2 (.ZN (XNOR_3_1_AND5_NUM2_OUT), .A1 (XNOR_1_3_AND5_NUM2_OUT), .A2 (GND));
      NOR2_X1 XNOR_3_2_AND5_NUM2 (.ZN (XNOR_3_2_AND5_NUM2_OUT), .A1 (GND), .A2 (XNOR_2_3_AND5_NUM2_OUT));
      NOR2_X1 XNOR_3_3_AND5_NUM2 (.ZN (XNOR_3_3_AND5_NUM2_OUT), .A1 (XNOR_3_1_AND5_NUM2_OUT), .A2 (XNOR_3_2_AND5_NUM2_OUT));

      wire XNOR_4_1_AND5_NUM2_OUT, XNOR_4_2_AND5_NUM2_OUT;
      NOR2_X1 XNOR_4_1_AND5_NUM2 (.ZN (XNOR_4_1_AND5_NUM2_OUT), .A1 (N986), .A2 (GND));
      NOR2_X1 XNOR_4_2_AND5_NUM2 (.ZN (XNOR_4_2_AND5_NUM2_OUT), .A1 (GND), .A2 (XNOR_3_3_AND5_NUM2_OUT));
      NOR2_X1 XNOR_4_3_AND5_NUM2 (.ZN (N1006), .A1 (XNOR_4_1_AND5_NUM2_OUT), .A2 (XNOR_4_2_AND5_NUM2_OUT));
      wire XNOR_1_1_AND5_NUM3_OUT, XNOR_1_2_AND5_NUM3_OUT, XNOR_1_3_AND5_NUM3_OUT;
      NOR2_X1 XNOR_1_1_AND5_NUM3 (.ZN (XNOR_1_1_AND5_NUM3_OUT), .A1 (N956), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND5_NUM3 (.ZN (XNOR_1_2_AND5_NUM3_OUT), .A1 (GND), .A2 (N886));
      NOR2_X1 XNOR_1_3_AND5_NUM3 (.ZN (XNOR_1_3_AND5_NUM3_OUT), .A1 (XNOR_1_1_AND5_NUM3_OUT), .A2 (XNOR_1_2_AND5_NUM3_OUT));

      wire XNOR_2_1_AND5_NUM3_OUT, XNOR_2_2_AND5_NUM3_OUT, XNOR_2_3_AND5_NUM3_OUT;
      NOR2_X1 XNOR_2_1_AND5_NUM3 (.ZN (XNOR_2_1_AND5_NUM3_OUT), .A1 (N957), .A2 (GND));
      NOR2_X1 XNOR_2_2_AND5_NUM3 (.ZN (XNOR_2_2_AND5_NUM3_OUT), .A1 (GND), .A2 (N899));
      NOR2_X1 XNOR_2_3_AND5_NUM3 (.ZN (XNOR_2_3_AND5_NUM3_OUT), .A1 (XNOR_2_1_AND5_NUM3_OUT), .A2 (XNOR_2_2_AND5_NUM3_OUT));

      wire XNOR_3_1_AND5_NUM3_OUT, XNOR_3_2_AND5_NUM3_OUT, XNOR_3_3_AND5_NUM3_OUT;
      NOR2_X1 XNOR_3_1_AND5_NUM3 (.ZN (XNOR_3_1_AND5_NUM3_OUT), .A1 (XNOR_1_3_AND5_NUM3_OUT), .A2 (GND));
      NOR2_X1 XNOR_3_2_AND5_NUM3 (.ZN (XNOR_3_2_AND5_NUM3_OUT), .A1 (GND), .A2 (XNOR_2_3_AND5_NUM3_OUT));
      NOR2_X1 XNOR_3_3_AND5_NUM3 (.ZN (XNOR_3_3_AND5_NUM3_OUT), .A1 (XNOR_3_1_AND5_NUM3_OUT), .A2 (XNOR_3_2_AND5_NUM3_OUT));

      wire XNOR_4_1_AND5_NUM3_OUT, XNOR_4_2_AND5_NUM3_OUT;
      NOR2_X1 XNOR_4_1_AND5_NUM3 (.ZN (XNOR_4_1_AND5_NUM3_OUT), .A1 (N986), .A2 (GND));
      NOR2_X1 XNOR_4_2_AND5_NUM3 (.ZN (XNOR_4_2_AND5_NUM3_OUT), .A1 (GND), .A2 (XNOR_3_3_AND5_NUM3_OUT));
      NOR2_X1 XNOR_4_3_AND5_NUM3 (.ZN (N1011), .A1 (XNOR_4_1_AND5_NUM3_OUT), .A2 (XNOR_4_2_AND5_NUM3_OUT));
      wire XNOR_1_1_AND5_NUM4_OUT, XNOR_1_2_AND5_NUM4_OUT, XNOR_1_3_AND5_NUM4_OUT;
      NOR2_X1 XNOR_1_1_AND5_NUM4 (.ZN (XNOR_1_1_AND5_NUM4_OUT), .A1 (N834), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND5_NUM4 (.ZN (XNOR_1_2_AND5_NUM4_OUT), .A1 (GND), .A2 (N970));
      NOR2_X1 XNOR_1_3_AND5_NUM4 (.ZN (XNOR_1_3_AND5_NUM4_OUT), .A1 (XNOR_1_1_AND5_NUM4_OUT), .A2 (XNOR_1_2_AND5_NUM4_OUT));

      wire XNOR_2_1_AND5_NUM4_OUT, XNOR_2_2_AND5_NUM4_OUT, XNOR_2_3_AND5_NUM4_OUT;
      NOR2_X1 XNOR_2_1_AND5_NUM4 (.ZN (XNOR_2_1_AND5_NUM4_OUT), .A1 (N860), .A2 (GND));
      NOR2_X1 XNOR_2_2_AND5_NUM4 (.ZN (XNOR_2_2_AND5_NUM4_OUT), .A1 (GND), .A2 (N971));
      NOR2_X1 XNOR_2_3_AND5_NUM4 (.ZN (XNOR_2_3_AND5_NUM4_OUT), .A1 (XNOR_2_1_AND5_NUM4_OUT), .A2 (XNOR_2_2_AND5_NUM4_OUT));

      wire XNOR_3_1_AND5_NUM4_OUT, XNOR_3_2_AND5_NUM4_OUT, XNOR_3_3_AND5_NUM4_OUT;
      NOR2_X1 XNOR_3_1_AND5_NUM4 (.ZN (XNOR_3_1_AND5_NUM4_OUT), .A1 (XNOR_1_3_AND5_NUM4_OUT), .A2 (GND));
      NOR2_X1 XNOR_3_2_AND5_NUM4 (.ZN (XNOR_3_2_AND5_NUM4_OUT), .A1 (GND), .A2 (XNOR_2_3_AND5_NUM4_OUT));
      NOR2_X1 XNOR_3_3_AND5_NUM4 (.ZN (XNOR_3_3_AND5_NUM4_OUT), .A1 (XNOR_3_1_AND5_NUM4_OUT), .A2 (XNOR_3_2_AND5_NUM4_OUT));

      wire XNOR_4_1_AND5_NUM4_OUT, XNOR_4_2_AND5_NUM4_OUT;
      NOR2_X1 XNOR_4_1_AND5_NUM4 (.ZN (XNOR_4_1_AND5_NUM4_OUT), .A1 (N991), .A2 (GND));
      NOR2_X1 XNOR_4_2_AND5_NUM4 (.ZN (XNOR_4_2_AND5_NUM4_OUT), .A1 (GND), .A2 (XNOR_3_3_AND5_NUM4_OUT));
      NOR2_X1 XNOR_4_3_AND5_NUM4 (.ZN (N1016), .A1 (XNOR_4_1_AND5_NUM4_OUT), .A2 (XNOR_4_2_AND5_NUM4_OUT));
      wire XNOR_1_1_AND5_NUM5_OUT, XNOR_1_2_AND5_NUM5_OUT, XNOR_1_3_AND5_NUM5_OUT;
      NOR2_X1 XNOR_1_1_AND5_NUM5 (.ZN (XNOR_1_1_AND5_NUM5_OUT), .A1 (N834), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND5_NUM5 (.ZN (XNOR_1_2_AND5_NUM5_OUT), .A1 (GND), .A2 (N972));
      NOR2_X1 XNOR_1_3_AND5_NUM5 (.ZN (XNOR_1_3_AND5_NUM5_OUT), .A1 (XNOR_1_1_AND5_NUM5_OUT), .A2 (XNOR_1_2_AND5_NUM5_OUT));

      wire XNOR_2_1_AND5_NUM5_OUT, XNOR_2_2_AND5_NUM5_OUT, XNOR_2_3_AND5_NUM5_OUT;
      NOR2_X1 XNOR_2_1_AND5_NUM5 (.ZN (XNOR_2_1_AND5_NUM5_OUT), .A1 (N973), .A2 (GND));
      NOR2_X1 XNOR_2_2_AND5_NUM5 (.ZN (XNOR_2_2_AND5_NUM5_OUT), .A1 (GND), .A2 (N873));
      NOR2_X1 XNOR_2_3_AND5_NUM5 (.ZN (XNOR_2_3_AND5_NUM5_OUT), .A1 (XNOR_2_1_AND5_NUM5_OUT), .A2 (XNOR_2_2_AND5_NUM5_OUT));

      wire XNOR_3_1_AND5_NUM5_OUT, XNOR_3_2_AND5_NUM5_OUT, XNOR_3_3_AND5_NUM5_OUT;
      NOR2_X1 XNOR_3_1_AND5_NUM5 (.ZN (XNOR_3_1_AND5_NUM5_OUT), .A1 (XNOR_1_3_AND5_NUM5_OUT), .A2 (GND));
      NOR2_X1 XNOR_3_2_AND5_NUM5 (.ZN (XNOR_3_2_AND5_NUM5_OUT), .A1 (GND), .A2 (XNOR_2_3_AND5_NUM5_OUT));
      NOR2_X1 XNOR_3_3_AND5_NUM5 (.ZN (XNOR_3_3_AND5_NUM5_OUT), .A1 (XNOR_3_1_AND5_NUM5_OUT), .A2 (XNOR_3_2_AND5_NUM5_OUT));

      wire XNOR_4_1_AND5_NUM5_OUT, XNOR_4_2_AND5_NUM5_OUT;
      NOR2_X1 XNOR_4_1_AND5_NUM5 (.ZN (XNOR_4_1_AND5_NUM5_OUT), .A1 (N991), .A2 (GND));
      NOR2_X1 XNOR_4_2_AND5_NUM5 (.ZN (XNOR_4_2_AND5_NUM5_OUT), .A1 (GND), .A2 (XNOR_3_3_AND5_NUM5_OUT));
      NOR2_X1 XNOR_4_3_AND5_NUM5 (.ZN (N1021), .A1 (XNOR_4_1_AND5_NUM5_OUT), .A2 (XNOR_4_2_AND5_NUM5_OUT));
      wire XNOR_1_1_AND5_NUM6_OUT, XNOR_1_2_AND5_NUM6_OUT, XNOR_1_3_AND5_NUM6_OUT;
      NOR2_X1 XNOR_1_1_AND5_NUM6 (.ZN (XNOR_1_1_AND5_NUM6_OUT), .A1 (N974), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND5_NUM6 (.ZN (XNOR_1_2_AND5_NUM6_OUT), .A1 (GND), .A2 (N847));
      NOR2_X1 XNOR_1_3_AND5_NUM6 (.ZN (XNOR_1_3_AND5_NUM6_OUT), .A1 (XNOR_1_1_AND5_NUM6_OUT), .A2 (XNOR_1_2_AND5_NUM6_OUT));

      wire XNOR_2_1_AND5_NUM6_OUT, XNOR_2_2_AND5_NUM6_OUT, XNOR_2_3_AND5_NUM6_OUT;
      NOR2_X1 XNOR_2_1_AND5_NUM6 (.ZN (XNOR_2_1_AND5_NUM6_OUT), .A1 (N860), .A2 (GND));
      NOR2_X1 XNOR_2_2_AND5_NUM6 (.ZN (XNOR_2_2_AND5_NUM6_OUT), .A1 (GND), .A2 (N975));
      NOR2_X1 XNOR_2_3_AND5_NUM6 (.ZN (XNOR_2_3_AND5_NUM6_OUT), .A1 (XNOR_2_1_AND5_NUM6_OUT), .A2 (XNOR_2_2_AND5_NUM6_OUT));

      wire XNOR_3_1_AND5_NUM6_OUT, XNOR_3_2_AND5_NUM6_OUT, XNOR_3_3_AND5_NUM6_OUT;
      NOR2_X1 XNOR_3_1_AND5_NUM6 (.ZN (XNOR_3_1_AND5_NUM6_OUT), .A1 (XNOR_1_3_AND5_NUM6_OUT), .A2 (GND));
      NOR2_X1 XNOR_3_2_AND5_NUM6 (.ZN (XNOR_3_2_AND5_NUM6_OUT), .A1 (GND), .A2 (XNOR_2_3_AND5_NUM6_OUT));
      NOR2_X1 XNOR_3_3_AND5_NUM6 (.ZN (XNOR_3_3_AND5_NUM6_OUT), .A1 (XNOR_3_1_AND5_NUM6_OUT), .A2 (XNOR_3_2_AND5_NUM6_OUT));

      wire XNOR_4_1_AND5_NUM6_OUT, XNOR_4_2_AND5_NUM6_OUT;
      NOR2_X1 XNOR_4_1_AND5_NUM6 (.ZN (XNOR_4_1_AND5_NUM6_OUT), .A1 (N991), .A2 (GND));
      NOR2_X1 XNOR_4_2_AND5_NUM6 (.ZN (XNOR_4_2_AND5_NUM6_OUT), .A1 (GND), .A2 (XNOR_3_3_AND5_NUM6_OUT));
      NOR2_X1 XNOR_4_3_AND5_NUM6 (.ZN (N1026), .A1 (XNOR_4_1_AND5_NUM6_OUT), .A2 (XNOR_4_2_AND5_NUM6_OUT));
      wire XNOR_1_1_AND5_NUM7_OUT, XNOR_1_2_AND5_NUM7_OUT, XNOR_1_3_AND5_NUM7_OUT;
      NOR2_X1 XNOR_1_1_AND5_NUM7 (.ZN (XNOR_1_1_AND5_NUM7_OUT), .A1 (N976), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND5_NUM7 (.ZN (XNOR_1_2_AND5_NUM7_OUT), .A1 (GND), .A2 (N847));
      NOR2_X1 XNOR_1_3_AND5_NUM7 (.ZN (XNOR_1_3_AND5_NUM7_OUT), .A1 (XNOR_1_1_AND5_NUM7_OUT), .A2 (XNOR_1_2_AND5_NUM7_OUT));

      wire XNOR_2_1_AND5_NUM7_OUT, XNOR_2_2_AND5_NUM7_OUT, XNOR_2_3_AND5_NUM7_OUT;
      NOR2_X1 XNOR_2_1_AND5_NUM7 (.ZN (XNOR_2_1_AND5_NUM7_OUT), .A1 (N977), .A2 (GND));
      NOR2_X1 XNOR_2_2_AND5_NUM7 (.ZN (XNOR_2_2_AND5_NUM7_OUT), .A1 (GND), .A2 (N873));
      NOR2_X1 XNOR_2_3_AND5_NUM7 (.ZN (XNOR_2_3_AND5_NUM7_OUT), .A1 (XNOR_2_1_AND5_NUM7_OUT), .A2 (XNOR_2_2_AND5_NUM7_OUT));

      wire XNOR_3_1_AND5_NUM7_OUT, XNOR_3_2_AND5_NUM7_OUT, XNOR_3_3_AND5_NUM7_OUT;
      NOR2_X1 XNOR_3_1_AND5_NUM7 (.ZN (XNOR_3_1_AND5_NUM7_OUT), .A1 (XNOR_1_3_AND5_NUM7_OUT), .A2 (GND));
      NOR2_X1 XNOR_3_2_AND5_NUM7 (.ZN (XNOR_3_2_AND5_NUM7_OUT), .A1 (GND), .A2 (XNOR_2_3_AND5_NUM7_OUT));
      NOR2_X1 XNOR_3_3_AND5_NUM7 (.ZN (XNOR_3_3_AND5_NUM7_OUT), .A1 (XNOR_3_1_AND5_NUM7_OUT), .A2 (XNOR_3_2_AND5_NUM7_OUT));

      wire XNOR_4_1_AND5_NUM7_OUT, XNOR_4_2_AND5_NUM7_OUT;
      NOR2_X1 XNOR_4_1_AND5_NUM7 (.ZN (XNOR_4_1_AND5_NUM7_OUT), .A1 (N991), .A2 (GND));
      NOR2_X1 XNOR_4_2_AND5_NUM7 (.ZN (XNOR_4_2_AND5_NUM7_OUT), .A1 (GND), .A2 (XNOR_3_3_AND5_NUM7_OUT));
      NOR2_X1 XNOR_4_3_AND5_NUM7 (.ZN (N1031), .A1 (XNOR_4_1_AND5_NUM7_OUT), .A2 (XNOR_4_2_AND5_NUM7_OUT));
      wire XNOR_1_1_AND2_NUM8_OUT, XNOR_1_2_AND2_NUM8_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM8 (.ZN (XNOR_1_1_AND2_NUM8_OUT), .A1 (N834), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM8 (.ZN (XNOR_1_2_AND2_NUM8_OUT), .A1 (GND), .A2 (N996));
      NOR2_X1 XNOR_1_3_AND2_NUM8 (.ZN (N1036), .A1 (XNOR_1_1_AND2_NUM8_OUT), .A2 (XNOR_1_2_AND2_NUM8_OUT));
      wire XNOR_1_1_AND2_NUM9_OUT, XNOR_1_2_AND2_NUM9_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM9 (.ZN (XNOR_1_1_AND2_NUM9_OUT), .A1 (N847), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM9 (.ZN (XNOR_1_2_AND2_NUM9_OUT), .A1 (GND), .A2 (N996));
      NOR2_X1 XNOR_1_3_AND2_NUM9 (.ZN (N1039), .A1 (XNOR_1_1_AND2_NUM9_OUT), .A2 (XNOR_1_2_AND2_NUM9_OUT));
      wire XNOR_1_1_AND2_NUM10_OUT, XNOR_1_2_AND2_NUM10_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM10 (.ZN (XNOR_1_1_AND2_NUM10_OUT), .A1 (N860), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM10 (.ZN (XNOR_1_2_AND2_NUM10_OUT), .A1 (GND), .A2 (N996));
      NOR2_X1 XNOR_1_3_AND2_NUM10 (.ZN (N1042), .A1 (XNOR_1_1_AND2_NUM10_OUT), .A2 (XNOR_1_2_AND2_NUM10_OUT));
      wire XNOR_1_1_AND2_NUM11_OUT, XNOR_1_2_AND2_NUM11_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM11 (.ZN (XNOR_1_1_AND2_NUM11_OUT), .A1 (N873), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM11 (.ZN (XNOR_1_2_AND2_NUM11_OUT), .A1 (GND), .A2 (N996));
      NOR2_X1 XNOR_1_3_AND2_NUM11 (.ZN (N1045), .A1 (XNOR_1_1_AND2_NUM11_OUT), .A2 (XNOR_1_2_AND2_NUM11_OUT));
      wire XNOR_1_1_AND2_NUM12_OUT, XNOR_1_2_AND2_NUM12_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM12 (.ZN (XNOR_1_1_AND2_NUM12_OUT), .A1 (N834), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM12 (.ZN (XNOR_1_2_AND2_NUM12_OUT), .A1 (GND), .A2 (N1001));
      NOR2_X1 XNOR_1_3_AND2_NUM12 (.ZN (N1048), .A1 (XNOR_1_1_AND2_NUM12_OUT), .A2 (XNOR_1_2_AND2_NUM12_OUT));
      wire XNOR_1_1_AND2_NUM13_OUT, XNOR_1_2_AND2_NUM13_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM13 (.ZN (XNOR_1_1_AND2_NUM13_OUT), .A1 (N847), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM13 (.ZN (XNOR_1_2_AND2_NUM13_OUT), .A1 (GND), .A2 (N1001));
      NOR2_X1 XNOR_1_3_AND2_NUM13 (.ZN (N1051), .A1 (XNOR_1_1_AND2_NUM13_OUT), .A2 (XNOR_1_2_AND2_NUM13_OUT));
      wire XNOR_1_1_AND2_NUM14_OUT, XNOR_1_2_AND2_NUM14_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM14 (.ZN (XNOR_1_1_AND2_NUM14_OUT), .A1 (N860), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM14 (.ZN (XNOR_1_2_AND2_NUM14_OUT), .A1 (GND), .A2 (N1001));
      NOR2_X1 XNOR_1_3_AND2_NUM14 (.ZN (N1054), .A1 (XNOR_1_1_AND2_NUM14_OUT), .A2 (XNOR_1_2_AND2_NUM14_OUT));
      wire XNOR_1_1_AND2_NUM15_OUT, XNOR_1_2_AND2_NUM15_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM15 (.ZN (XNOR_1_1_AND2_NUM15_OUT), .A1 (N873), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM15 (.ZN (XNOR_1_2_AND2_NUM15_OUT), .A1 (GND), .A2 (N1001));
      NOR2_X1 XNOR_1_3_AND2_NUM15 (.ZN (N1057), .A1 (XNOR_1_1_AND2_NUM15_OUT), .A2 (XNOR_1_2_AND2_NUM15_OUT));
      wire XNOR_1_1_AND2_NUM16_OUT, XNOR_1_2_AND2_NUM16_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM16 (.ZN (XNOR_1_1_AND2_NUM16_OUT), .A1 (N834), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM16 (.ZN (XNOR_1_2_AND2_NUM16_OUT), .A1 (GND), .A2 (N1006));
      NOR2_X1 XNOR_1_3_AND2_NUM16 (.ZN (N1060), .A1 (XNOR_1_1_AND2_NUM16_OUT), .A2 (XNOR_1_2_AND2_NUM16_OUT));
      wire XNOR_1_1_AND2_NUM17_OUT, XNOR_1_2_AND2_NUM17_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM17 (.ZN (XNOR_1_1_AND2_NUM17_OUT), .A1 (N847), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM17 (.ZN (XNOR_1_2_AND2_NUM17_OUT), .A1 (GND), .A2 (N1006));
      NOR2_X1 XNOR_1_3_AND2_NUM17 (.ZN (N1063), .A1 (XNOR_1_1_AND2_NUM17_OUT), .A2 (XNOR_1_2_AND2_NUM17_OUT));
      wire XNOR_1_1_AND2_NUM18_OUT, XNOR_1_2_AND2_NUM18_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM18 (.ZN (XNOR_1_1_AND2_NUM18_OUT), .A1 (N860), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM18 (.ZN (XNOR_1_2_AND2_NUM18_OUT), .A1 (GND), .A2 (N1006));
      NOR2_X1 XNOR_1_3_AND2_NUM18 (.ZN (N1066), .A1 (XNOR_1_1_AND2_NUM18_OUT), .A2 (XNOR_1_2_AND2_NUM18_OUT));
      wire XNOR_1_1_AND2_NUM19_OUT, XNOR_1_2_AND2_NUM19_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM19 (.ZN (XNOR_1_1_AND2_NUM19_OUT), .A1 (N873), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM19 (.ZN (XNOR_1_2_AND2_NUM19_OUT), .A1 (GND), .A2 (N1006));
      NOR2_X1 XNOR_1_3_AND2_NUM19 (.ZN (N1069), .A1 (XNOR_1_1_AND2_NUM19_OUT), .A2 (XNOR_1_2_AND2_NUM19_OUT));
      wire XNOR_1_1_AND2_NUM20_OUT, XNOR_1_2_AND2_NUM20_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM20 (.ZN (XNOR_1_1_AND2_NUM20_OUT), .A1 (N834), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM20 (.ZN (XNOR_1_2_AND2_NUM20_OUT), .A1 (GND), .A2 (N1011));
      NOR2_X1 XNOR_1_3_AND2_NUM20 (.ZN (N1072), .A1 (XNOR_1_1_AND2_NUM20_OUT), .A2 (XNOR_1_2_AND2_NUM20_OUT));
      wire XNOR_1_1_AND2_NUM21_OUT, XNOR_1_2_AND2_NUM21_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM21 (.ZN (XNOR_1_1_AND2_NUM21_OUT), .A1 (N847), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM21 (.ZN (XNOR_1_2_AND2_NUM21_OUT), .A1 (GND), .A2 (N1011));
      NOR2_X1 XNOR_1_3_AND2_NUM21 (.ZN (N1075), .A1 (XNOR_1_1_AND2_NUM21_OUT), .A2 (XNOR_1_2_AND2_NUM21_OUT));
      wire XNOR_1_1_AND2_NUM22_OUT, XNOR_1_2_AND2_NUM22_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM22 (.ZN (XNOR_1_1_AND2_NUM22_OUT), .A1 (N860), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM22 (.ZN (XNOR_1_2_AND2_NUM22_OUT), .A1 (GND), .A2 (N1011));
      NOR2_X1 XNOR_1_3_AND2_NUM22 (.ZN (N1078), .A1 (XNOR_1_1_AND2_NUM22_OUT), .A2 (XNOR_1_2_AND2_NUM22_OUT));
      wire XNOR_1_1_AND2_NUM23_OUT, XNOR_1_2_AND2_NUM23_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM23 (.ZN (XNOR_1_1_AND2_NUM23_OUT), .A1 (N873), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM23 (.ZN (XNOR_1_2_AND2_NUM23_OUT), .A1 (GND), .A2 (N1011));
      NOR2_X1 XNOR_1_3_AND2_NUM23 (.ZN (N1081), .A1 (XNOR_1_1_AND2_NUM23_OUT), .A2 (XNOR_1_2_AND2_NUM23_OUT));
      wire XNOR_1_1_AND2_NUM24_OUT, XNOR_1_2_AND2_NUM24_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM24 (.ZN (XNOR_1_1_AND2_NUM24_OUT), .A1 (N925), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM24 (.ZN (XNOR_1_2_AND2_NUM24_OUT), .A1 (GND), .A2 (N1016));
      NOR2_X1 XNOR_1_3_AND2_NUM24 (.ZN (N1084), .A1 (XNOR_1_1_AND2_NUM24_OUT), .A2 (XNOR_1_2_AND2_NUM24_OUT));
      wire XNOR_1_1_AND2_NUM25_OUT, XNOR_1_2_AND2_NUM25_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM25 (.ZN (XNOR_1_1_AND2_NUM25_OUT), .A1 (N886), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM25 (.ZN (XNOR_1_2_AND2_NUM25_OUT), .A1 (GND), .A2 (N1016));
      NOR2_X1 XNOR_1_3_AND2_NUM25 (.ZN (N1087), .A1 (XNOR_1_1_AND2_NUM25_OUT), .A2 (XNOR_1_2_AND2_NUM25_OUT));
      wire XNOR_1_1_AND2_NUM26_OUT, XNOR_1_2_AND2_NUM26_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM26 (.ZN (XNOR_1_1_AND2_NUM26_OUT), .A1 (N912), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM26 (.ZN (XNOR_1_2_AND2_NUM26_OUT), .A1 (GND), .A2 (N1016));
      NOR2_X1 XNOR_1_3_AND2_NUM26 (.ZN (N1090), .A1 (XNOR_1_1_AND2_NUM26_OUT), .A2 (XNOR_1_2_AND2_NUM26_OUT));
      wire XNOR_1_1_AND2_NUM27_OUT, XNOR_1_2_AND2_NUM27_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM27 (.ZN (XNOR_1_1_AND2_NUM27_OUT), .A1 (N899), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM27 (.ZN (XNOR_1_2_AND2_NUM27_OUT), .A1 (GND), .A2 (N1016));
      NOR2_X1 XNOR_1_3_AND2_NUM27 (.ZN (N1093), .A1 (XNOR_1_1_AND2_NUM27_OUT), .A2 (XNOR_1_2_AND2_NUM27_OUT));
      wire XNOR_1_1_AND2_NUM28_OUT, XNOR_1_2_AND2_NUM28_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM28 (.ZN (XNOR_1_1_AND2_NUM28_OUT), .A1 (N925), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM28 (.ZN (XNOR_1_2_AND2_NUM28_OUT), .A1 (GND), .A2 (N1021));
      NOR2_X1 XNOR_1_3_AND2_NUM28 (.ZN (N1096), .A1 (XNOR_1_1_AND2_NUM28_OUT), .A2 (XNOR_1_2_AND2_NUM28_OUT));
      wire XNOR_1_1_AND2_NUM29_OUT, XNOR_1_2_AND2_NUM29_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM29 (.ZN (XNOR_1_1_AND2_NUM29_OUT), .A1 (N886), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM29 (.ZN (XNOR_1_2_AND2_NUM29_OUT), .A1 (GND), .A2 (N1021));
      NOR2_X1 XNOR_1_3_AND2_NUM29 (.ZN (N1099), .A1 (XNOR_1_1_AND2_NUM29_OUT), .A2 (XNOR_1_2_AND2_NUM29_OUT));
      wire XNOR_1_1_AND2_NUM30_OUT, XNOR_1_2_AND2_NUM30_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM30 (.ZN (XNOR_1_1_AND2_NUM30_OUT), .A1 (N912), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM30 (.ZN (XNOR_1_2_AND2_NUM30_OUT), .A1 (GND), .A2 (N1021));
      NOR2_X1 XNOR_1_3_AND2_NUM30 (.ZN (N1102), .A1 (XNOR_1_1_AND2_NUM30_OUT), .A2 (XNOR_1_2_AND2_NUM30_OUT));
      wire XNOR_1_1_AND2_NUM31_OUT, XNOR_1_2_AND2_NUM31_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM31 (.ZN (XNOR_1_1_AND2_NUM31_OUT), .A1 (N899), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM31 (.ZN (XNOR_1_2_AND2_NUM31_OUT), .A1 (GND), .A2 (N1021));
      NOR2_X1 XNOR_1_3_AND2_NUM31 (.ZN (N1105), .A1 (XNOR_1_1_AND2_NUM31_OUT), .A2 (XNOR_1_2_AND2_NUM31_OUT));
      wire XNOR_1_1_AND2_NUM32_OUT, XNOR_1_2_AND2_NUM32_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM32 (.ZN (XNOR_1_1_AND2_NUM32_OUT), .A1 (N925), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM32 (.ZN (XNOR_1_2_AND2_NUM32_OUT), .A1 (GND), .A2 (N1026));
      NOR2_X1 XNOR_1_3_AND2_NUM32 (.ZN (N1108), .A1 (XNOR_1_1_AND2_NUM32_OUT), .A2 (XNOR_1_2_AND2_NUM32_OUT));
      wire XNOR_1_1_AND2_NUM33_OUT, XNOR_1_2_AND2_NUM33_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM33 (.ZN (XNOR_1_1_AND2_NUM33_OUT), .A1 (N886), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM33 (.ZN (XNOR_1_2_AND2_NUM33_OUT), .A1 (GND), .A2 (N1026));
      NOR2_X1 XNOR_1_3_AND2_NUM33 (.ZN (N1111), .A1 (XNOR_1_1_AND2_NUM33_OUT), .A2 (XNOR_1_2_AND2_NUM33_OUT));
      wire XNOR_1_1_AND2_NUM34_OUT, XNOR_1_2_AND2_NUM34_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM34 (.ZN (XNOR_1_1_AND2_NUM34_OUT), .A1 (N912), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM34 (.ZN (XNOR_1_2_AND2_NUM34_OUT), .A1 (GND), .A2 (N1026));
      NOR2_X1 XNOR_1_3_AND2_NUM34 (.ZN (N1114), .A1 (XNOR_1_1_AND2_NUM34_OUT), .A2 (XNOR_1_2_AND2_NUM34_OUT));
      wire XNOR_1_1_AND2_NUM35_OUT, XNOR_1_2_AND2_NUM35_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM35 (.ZN (XNOR_1_1_AND2_NUM35_OUT), .A1 (N899), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM35 (.ZN (XNOR_1_2_AND2_NUM35_OUT), .A1 (GND), .A2 (N1026));
      NOR2_X1 XNOR_1_3_AND2_NUM35 (.ZN (N1117), .A1 (XNOR_1_1_AND2_NUM35_OUT), .A2 (XNOR_1_2_AND2_NUM35_OUT));
      wire XNOR_1_1_AND2_NUM36_OUT, XNOR_1_2_AND2_NUM36_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM36 (.ZN (XNOR_1_1_AND2_NUM36_OUT), .A1 (N925), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM36 (.ZN (XNOR_1_2_AND2_NUM36_OUT), .A1 (GND), .A2 (N1031));
      NOR2_X1 XNOR_1_3_AND2_NUM36 (.ZN (N1120), .A1 (XNOR_1_1_AND2_NUM36_OUT), .A2 (XNOR_1_2_AND2_NUM36_OUT));
      wire XNOR_1_1_AND2_NUM37_OUT, XNOR_1_2_AND2_NUM37_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM37 (.ZN (XNOR_1_1_AND2_NUM37_OUT), .A1 (N886), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM37 (.ZN (XNOR_1_2_AND2_NUM37_OUT), .A1 (GND), .A2 (N1031));
      NOR2_X1 XNOR_1_3_AND2_NUM37 (.ZN (N1123), .A1 (XNOR_1_1_AND2_NUM37_OUT), .A2 (XNOR_1_2_AND2_NUM37_OUT));
      wire XNOR_1_1_AND2_NUM38_OUT, XNOR_1_2_AND2_NUM38_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM38 (.ZN (XNOR_1_1_AND2_NUM38_OUT), .A1 (N912), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM38 (.ZN (XNOR_1_2_AND2_NUM38_OUT), .A1 (GND), .A2 (N1031));
      NOR2_X1 XNOR_1_3_AND2_NUM38 (.ZN (N1126), .A1 (XNOR_1_1_AND2_NUM38_OUT), .A2 (XNOR_1_2_AND2_NUM38_OUT));
      wire XNOR_1_1_AND2_NUM39_OUT, XNOR_1_2_AND2_NUM39_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM39 (.ZN (XNOR_1_1_AND2_NUM39_OUT), .A1 (N899), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM39 (.ZN (XNOR_1_2_AND2_NUM39_OUT), .A1 (GND), .A2 (N1031));
      NOR2_X1 XNOR_1_3_AND2_NUM39 (.ZN (N1129), .A1 (XNOR_1_1_AND2_NUM39_OUT), .A2 (XNOR_1_2_AND2_NUM39_OUT));
      wire XNOR_1_1_NAND2_NUM288_OUT, XNOR_1_2_NAND2_NUM288_OUT, XNOR_1_3_NAND2_NUM288_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM288 (.ZN (XNOR_1_1_NAND2_NUM288_OUT), .A1 (N1), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM288 (.ZN (XNOR_1_2_NAND2_NUM288_OUT), .A1 (GND), .A2 (N1036));
      NOR2_X1 XNOR_1_3_NAND2_NUM288 (.ZN (XNOR_1_3_NAND2_NUM288_OUT), .A1 (XNOR_1_1_NAND2_NUM288_OUT), .A2 (XNOR_1_2_NAND2_NUM288_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM288 (.ZN (N1132), .A1 (XNOR_1_3_NAND2_NUM288_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM289_OUT, XNOR_1_2_NAND2_NUM289_OUT, XNOR_1_3_NAND2_NUM289_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM289 (.ZN (XNOR_1_1_NAND2_NUM289_OUT), .A1 (N8), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM289 (.ZN (XNOR_1_2_NAND2_NUM289_OUT), .A1 (GND), .A2 (N1039));
      NOR2_X1 XNOR_1_3_NAND2_NUM289 (.ZN (XNOR_1_3_NAND2_NUM289_OUT), .A1 (XNOR_1_1_NAND2_NUM289_OUT), .A2 (XNOR_1_2_NAND2_NUM289_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM289 (.ZN (N1135), .A1 (XNOR_1_3_NAND2_NUM289_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM290_OUT, XNOR_1_2_NAND2_NUM290_OUT, XNOR_1_3_NAND2_NUM290_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM290 (.ZN (XNOR_1_1_NAND2_NUM290_OUT), .A1 (N15), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM290 (.ZN (XNOR_1_2_NAND2_NUM290_OUT), .A1 (GND), .A2 (N1042));
      NOR2_X1 XNOR_1_3_NAND2_NUM290 (.ZN (XNOR_1_3_NAND2_NUM290_OUT), .A1 (XNOR_1_1_NAND2_NUM290_OUT), .A2 (XNOR_1_2_NAND2_NUM290_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM290 (.ZN (N1138), .A1 (XNOR_1_3_NAND2_NUM290_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM291_OUT, XNOR_1_2_NAND2_NUM291_OUT, XNOR_1_3_NAND2_NUM291_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM291 (.ZN (XNOR_1_1_NAND2_NUM291_OUT), .A1 (N22), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM291 (.ZN (XNOR_1_2_NAND2_NUM291_OUT), .A1 (GND), .A2 (N1045));
      NOR2_X1 XNOR_1_3_NAND2_NUM291 (.ZN (XNOR_1_3_NAND2_NUM291_OUT), .A1 (XNOR_1_1_NAND2_NUM291_OUT), .A2 (XNOR_1_2_NAND2_NUM291_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM291 (.ZN (N1141), .A1 (XNOR_1_3_NAND2_NUM291_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM292_OUT, XNOR_1_2_NAND2_NUM292_OUT, XNOR_1_3_NAND2_NUM292_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM292 (.ZN (XNOR_1_1_NAND2_NUM292_OUT), .A1 (N29), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM292 (.ZN (XNOR_1_2_NAND2_NUM292_OUT), .A1 (GND), .A2 (N1048));
      NOR2_X1 XNOR_1_3_NAND2_NUM292 (.ZN (XNOR_1_3_NAND2_NUM292_OUT), .A1 (XNOR_1_1_NAND2_NUM292_OUT), .A2 (XNOR_1_2_NAND2_NUM292_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM292 (.ZN (N1144), .A1 (XNOR_1_3_NAND2_NUM292_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM293_OUT, XNOR_1_2_NAND2_NUM293_OUT, XNOR_1_3_NAND2_NUM293_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM293 (.ZN (XNOR_1_1_NAND2_NUM293_OUT), .A1 (N36), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM293 (.ZN (XNOR_1_2_NAND2_NUM293_OUT), .A1 (GND), .A2 (N1051));
      NOR2_X1 XNOR_1_3_NAND2_NUM293 (.ZN (XNOR_1_3_NAND2_NUM293_OUT), .A1 (XNOR_1_1_NAND2_NUM293_OUT), .A2 (XNOR_1_2_NAND2_NUM293_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM293 (.ZN (N1147), .A1 (XNOR_1_3_NAND2_NUM293_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM294_OUT, XNOR_1_2_NAND2_NUM294_OUT, XNOR_1_3_NAND2_NUM294_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM294 (.ZN (XNOR_1_1_NAND2_NUM294_OUT), .A1 (N43), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM294 (.ZN (XNOR_1_2_NAND2_NUM294_OUT), .A1 (GND), .A2 (N1054));
      NOR2_X1 XNOR_1_3_NAND2_NUM294 (.ZN (XNOR_1_3_NAND2_NUM294_OUT), .A1 (XNOR_1_1_NAND2_NUM294_OUT), .A2 (XNOR_1_2_NAND2_NUM294_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM294 (.ZN (N1150), .A1 (XNOR_1_3_NAND2_NUM294_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM295_OUT, XNOR_1_2_NAND2_NUM295_OUT, XNOR_1_3_NAND2_NUM295_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM295 (.ZN (XNOR_1_1_NAND2_NUM295_OUT), .A1 (N50), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM295 (.ZN (XNOR_1_2_NAND2_NUM295_OUT), .A1 (GND), .A2 (N1057));
      NOR2_X1 XNOR_1_3_NAND2_NUM295 (.ZN (XNOR_1_3_NAND2_NUM295_OUT), .A1 (XNOR_1_1_NAND2_NUM295_OUT), .A2 (XNOR_1_2_NAND2_NUM295_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM295 (.ZN (N1153), .A1 (XNOR_1_3_NAND2_NUM295_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM296_OUT, XNOR_1_2_NAND2_NUM296_OUT, XNOR_1_3_NAND2_NUM296_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM296 (.ZN (XNOR_1_1_NAND2_NUM296_OUT), .A1 (N57), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM296 (.ZN (XNOR_1_2_NAND2_NUM296_OUT), .A1 (GND), .A2 (N1060));
      NOR2_X1 XNOR_1_3_NAND2_NUM296 (.ZN (XNOR_1_3_NAND2_NUM296_OUT), .A1 (XNOR_1_1_NAND2_NUM296_OUT), .A2 (XNOR_1_2_NAND2_NUM296_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM296 (.ZN (N1156), .A1 (XNOR_1_3_NAND2_NUM296_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM297_OUT, XNOR_1_2_NAND2_NUM297_OUT, XNOR_1_3_NAND2_NUM297_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM297 (.ZN (XNOR_1_1_NAND2_NUM297_OUT), .A1 (N64), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM297 (.ZN (XNOR_1_2_NAND2_NUM297_OUT), .A1 (GND), .A2 (N1063));
      NOR2_X1 XNOR_1_3_NAND2_NUM297 (.ZN (XNOR_1_3_NAND2_NUM297_OUT), .A1 (XNOR_1_1_NAND2_NUM297_OUT), .A2 (XNOR_1_2_NAND2_NUM297_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM297 (.ZN (N1159), .A1 (XNOR_1_3_NAND2_NUM297_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM298_OUT, XNOR_1_2_NAND2_NUM298_OUT, XNOR_1_3_NAND2_NUM298_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM298 (.ZN (XNOR_1_1_NAND2_NUM298_OUT), .A1 (N71), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM298 (.ZN (XNOR_1_2_NAND2_NUM298_OUT), .A1 (GND), .A2 (N1066));
      NOR2_X1 XNOR_1_3_NAND2_NUM298 (.ZN (XNOR_1_3_NAND2_NUM298_OUT), .A1 (XNOR_1_1_NAND2_NUM298_OUT), .A2 (XNOR_1_2_NAND2_NUM298_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM298 (.ZN (N1162), .A1 (XNOR_1_3_NAND2_NUM298_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM299_OUT, XNOR_1_2_NAND2_NUM299_OUT, XNOR_1_3_NAND2_NUM299_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM299 (.ZN (XNOR_1_1_NAND2_NUM299_OUT), .A1 (N78), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM299 (.ZN (XNOR_1_2_NAND2_NUM299_OUT), .A1 (GND), .A2 (N1069));
      NOR2_X1 XNOR_1_3_NAND2_NUM299 (.ZN (XNOR_1_3_NAND2_NUM299_OUT), .A1 (XNOR_1_1_NAND2_NUM299_OUT), .A2 (XNOR_1_2_NAND2_NUM299_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM299 (.ZN (N1165), .A1 (XNOR_1_3_NAND2_NUM299_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM300_OUT, XNOR_1_2_NAND2_NUM300_OUT, XNOR_1_3_NAND2_NUM300_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM300 (.ZN (XNOR_1_1_NAND2_NUM300_OUT), .A1 (N85), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM300 (.ZN (XNOR_1_2_NAND2_NUM300_OUT), .A1 (GND), .A2 (N1072));
      NOR2_X1 XNOR_1_3_NAND2_NUM300 (.ZN (XNOR_1_3_NAND2_NUM300_OUT), .A1 (XNOR_1_1_NAND2_NUM300_OUT), .A2 (XNOR_1_2_NAND2_NUM300_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM300 (.ZN (N1168), .A1 (XNOR_1_3_NAND2_NUM300_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM301_OUT, XNOR_1_2_NAND2_NUM301_OUT, XNOR_1_3_NAND2_NUM301_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM301 (.ZN (XNOR_1_1_NAND2_NUM301_OUT), .A1 (N92), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM301 (.ZN (XNOR_1_2_NAND2_NUM301_OUT), .A1 (GND), .A2 (N1075));
      NOR2_X1 XNOR_1_3_NAND2_NUM301 (.ZN (XNOR_1_3_NAND2_NUM301_OUT), .A1 (XNOR_1_1_NAND2_NUM301_OUT), .A2 (XNOR_1_2_NAND2_NUM301_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM301 (.ZN (N1171), .A1 (XNOR_1_3_NAND2_NUM301_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM302_OUT, XNOR_1_2_NAND2_NUM302_OUT, XNOR_1_3_NAND2_NUM302_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM302 (.ZN (XNOR_1_1_NAND2_NUM302_OUT), .A1 (N99), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM302 (.ZN (XNOR_1_2_NAND2_NUM302_OUT), .A1 (GND), .A2 (N1078));
      NOR2_X1 XNOR_1_3_NAND2_NUM302 (.ZN (XNOR_1_3_NAND2_NUM302_OUT), .A1 (XNOR_1_1_NAND2_NUM302_OUT), .A2 (XNOR_1_2_NAND2_NUM302_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM302 (.ZN (N1174), .A1 (XNOR_1_3_NAND2_NUM302_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM303_OUT, XNOR_1_2_NAND2_NUM303_OUT, XNOR_1_3_NAND2_NUM303_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM303 (.ZN (XNOR_1_1_NAND2_NUM303_OUT), .A1 (N106), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM303 (.ZN (XNOR_1_2_NAND2_NUM303_OUT), .A1 (GND), .A2 (N1081));
      NOR2_X1 XNOR_1_3_NAND2_NUM303 (.ZN (XNOR_1_3_NAND2_NUM303_OUT), .A1 (XNOR_1_1_NAND2_NUM303_OUT), .A2 (XNOR_1_2_NAND2_NUM303_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM303 (.ZN (N1177), .A1 (XNOR_1_3_NAND2_NUM303_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM304_OUT, XNOR_1_2_NAND2_NUM304_OUT, XNOR_1_3_NAND2_NUM304_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM304 (.ZN (XNOR_1_1_NAND2_NUM304_OUT), .A1 (N113), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM304 (.ZN (XNOR_1_2_NAND2_NUM304_OUT), .A1 (GND), .A2 (N1084));
      NOR2_X1 XNOR_1_3_NAND2_NUM304 (.ZN (XNOR_1_3_NAND2_NUM304_OUT), .A1 (XNOR_1_1_NAND2_NUM304_OUT), .A2 (XNOR_1_2_NAND2_NUM304_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM304 (.ZN (N1180), .A1 (XNOR_1_3_NAND2_NUM304_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM305_OUT, XNOR_1_2_NAND2_NUM305_OUT, XNOR_1_3_NAND2_NUM305_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM305 (.ZN (XNOR_1_1_NAND2_NUM305_OUT), .A1 (N120), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM305 (.ZN (XNOR_1_2_NAND2_NUM305_OUT), .A1 (GND), .A2 (N1087));
      NOR2_X1 XNOR_1_3_NAND2_NUM305 (.ZN (XNOR_1_3_NAND2_NUM305_OUT), .A1 (XNOR_1_1_NAND2_NUM305_OUT), .A2 (XNOR_1_2_NAND2_NUM305_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM305 (.ZN (N1183), .A1 (XNOR_1_3_NAND2_NUM305_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM306_OUT, XNOR_1_2_NAND2_NUM306_OUT, XNOR_1_3_NAND2_NUM306_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM306 (.ZN (XNOR_1_1_NAND2_NUM306_OUT), .A1 (N127), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM306 (.ZN (XNOR_1_2_NAND2_NUM306_OUT), .A1 (GND), .A2 (N1090));
      NOR2_X1 XNOR_1_3_NAND2_NUM306 (.ZN (XNOR_1_3_NAND2_NUM306_OUT), .A1 (XNOR_1_1_NAND2_NUM306_OUT), .A2 (XNOR_1_2_NAND2_NUM306_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM306 (.ZN (N1186), .A1 (XNOR_1_3_NAND2_NUM306_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM307_OUT, XNOR_1_2_NAND2_NUM307_OUT, XNOR_1_3_NAND2_NUM307_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM307 (.ZN (XNOR_1_1_NAND2_NUM307_OUT), .A1 (N134), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM307 (.ZN (XNOR_1_2_NAND2_NUM307_OUT), .A1 (GND), .A2 (N1093));
      NOR2_X1 XNOR_1_3_NAND2_NUM307 (.ZN (XNOR_1_3_NAND2_NUM307_OUT), .A1 (XNOR_1_1_NAND2_NUM307_OUT), .A2 (XNOR_1_2_NAND2_NUM307_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM307 (.ZN (N1189), .A1 (XNOR_1_3_NAND2_NUM307_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM308_OUT, XNOR_1_2_NAND2_NUM308_OUT, XNOR_1_3_NAND2_NUM308_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM308 (.ZN (XNOR_1_1_NAND2_NUM308_OUT), .A1 (N141), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM308 (.ZN (XNOR_1_2_NAND2_NUM308_OUT), .A1 (GND), .A2 (N1096));
      NOR2_X1 XNOR_1_3_NAND2_NUM308 (.ZN (XNOR_1_3_NAND2_NUM308_OUT), .A1 (XNOR_1_1_NAND2_NUM308_OUT), .A2 (XNOR_1_2_NAND2_NUM308_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM308 (.ZN (N1192), .A1 (XNOR_1_3_NAND2_NUM308_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM309_OUT, XNOR_1_2_NAND2_NUM309_OUT, XNOR_1_3_NAND2_NUM309_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM309 (.ZN (XNOR_1_1_NAND2_NUM309_OUT), .A1 (N148), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM309 (.ZN (XNOR_1_2_NAND2_NUM309_OUT), .A1 (GND), .A2 (N1099));
      NOR2_X1 XNOR_1_3_NAND2_NUM309 (.ZN (XNOR_1_3_NAND2_NUM309_OUT), .A1 (XNOR_1_1_NAND2_NUM309_OUT), .A2 (XNOR_1_2_NAND2_NUM309_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM309 (.ZN (N1195), .A1 (XNOR_1_3_NAND2_NUM309_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM310_OUT, XNOR_1_2_NAND2_NUM310_OUT, XNOR_1_3_NAND2_NUM310_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM310 (.ZN (XNOR_1_1_NAND2_NUM310_OUT), .A1 (N155), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM310 (.ZN (XNOR_1_2_NAND2_NUM310_OUT), .A1 (GND), .A2 (N1102));
      NOR2_X1 XNOR_1_3_NAND2_NUM310 (.ZN (XNOR_1_3_NAND2_NUM310_OUT), .A1 (XNOR_1_1_NAND2_NUM310_OUT), .A2 (XNOR_1_2_NAND2_NUM310_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM310 (.ZN (N1198), .A1 (XNOR_1_3_NAND2_NUM310_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM311_OUT, XNOR_1_2_NAND2_NUM311_OUT, XNOR_1_3_NAND2_NUM311_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM311 (.ZN (XNOR_1_1_NAND2_NUM311_OUT), .A1 (N162), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM311 (.ZN (XNOR_1_2_NAND2_NUM311_OUT), .A1 (GND), .A2 (N1105));
      NOR2_X1 XNOR_1_3_NAND2_NUM311 (.ZN (XNOR_1_3_NAND2_NUM311_OUT), .A1 (XNOR_1_1_NAND2_NUM311_OUT), .A2 (XNOR_1_2_NAND2_NUM311_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM311 (.ZN (N1201), .A1 (XNOR_1_3_NAND2_NUM311_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM312_OUT, XNOR_1_2_NAND2_NUM312_OUT, XNOR_1_3_NAND2_NUM312_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM312 (.ZN (XNOR_1_1_NAND2_NUM312_OUT), .A1 (N169), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM312 (.ZN (XNOR_1_2_NAND2_NUM312_OUT), .A1 (GND), .A2 (N1108));
      NOR2_X1 XNOR_1_3_NAND2_NUM312 (.ZN (XNOR_1_3_NAND2_NUM312_OUT), .A1 (XNOR_1_1_NAND2_NUM312_OUT), .A2 (XNOR_1_2_NAND2_NUM312_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM312 (.ZN (N1204), .A1 (XNOR_1_3_NAND2_NUM312_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM313_OUT, XNOR_1_2_NAND2_NUM313_OUT, XNOR_1_3_NAND2_NUM313_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM313 (.ZN (XNOR_1_1_NAND2_NUM313_OUT), .A1 (N176), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM313 (.ZN (XNOR_1_2_NAND2_NUM313_OUT), .A1 (GND), .A2 (N1111));
      NOR2_X1 XNOR_1_3_NAND2_NUM313 (.ZN (XNOR_1_3_NAND2_NUM313_OUT), .A1 (XNOR_1_1_NAND2_NUM313_OUT), .A2 (XNOR_1_2_NAND2_NUM313_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM313 (.ZN (N1207), .A1 (XNOR_1_3_NAND2_NUM313_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM314_OUT, XNOR_1_2_NAND2_NUM314_OUT, XNOR_1_3_NAND2_NUM314_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM314 (.ZN (XNOR_1_1_NAND2_NUM314_OUT), .A1 (N183), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM314 (.ZN (XNOR_1_2_NAND2_NUM314_OUT), .A1 (GND), .A2 (N1114));
      NOR2_X1 XNOR_1_3_NAND2_NUM314 (.ZN (XNOR_1_3_NAND2_NUM314_OUT), .A1 (XNOR_1_1_NAND2_NUM314_OUT), .A2 (XNOR_1_2_NAND2_NUM314_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM314 (.ZN (N1210), .A1 (XNOR_1_3_NAND2_NUM314_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM315_OUT, XNOR_1_2_NAND2_NUM315_OUT, XNOR_1_3_NAND2_NUM315_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM315 (.ZN (XNOR_1_1_NAND2_NUM315_OUT), .A1 (N190), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM315 (.ZN (XNOR_1_2_NAND2_NUM315_OUT), .A1 (GND), .A2 (N1117));
      NOR2_X1 XNOR_1_3_NAND2_NUM315 (.ZN (XNOR_1_3_NAND2_NUM315_OUT), .A1 (XNOR_1_1_NAND2_NUM315_OUT), .A2 (XNOR_1_2_NAND2_NUM315_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM315 (.ZN (N1213), .A1 (XNOR_1_3_NAND2_NUM315_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM316_OUT, XNOR_1_2_NAND2_NUM316_OUT, XNOR_1_3_NAND2_NUM316_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM316 (.ZN (XNOR_1_1_NAND2_NUM316_OUT), .A1 (N197), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM316 (.ZN (XNOR_1_2_NAND2_NUM316_OUT), .A1 (GND), .A2 (N1120));
      NOR2_X1 XNOR_1_3_NAND2_NUM316 (.ZN (XNOR_1_3_NAND2_NUM316_OUT), .A1 (XNOR_1_1_NAND2_NUM316_OUT), .A2 (XNOR_1_2_NAND2_NUM316_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM316 (.ZN (N1216), .A1 (XNOR_1_3_NAND2_NUM316_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM317_OUT, XNOR_1_2_NAND2_NUM317_OUT, XNOR_1_3_NAND2_NUM317_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM317 (.ZN (XNOR_1_1_NAND2_NUM317_OUT), .A1 (N204), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM317 (.ZN (XNOR_1_2_NAND2_NUM317_OUT), .A1 (GND), .A2 (N1123));
      NOR2_X1 XNOR_1_3_NAND2_NUM317 (.ZN (XNOR_1_3_NAND2_NUM317_OUT), .A1 (XNOR_1_1_NAND2_NUM317_OUT), .A2 (XNOR_1_2_NAND2_NUM317_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM317 (.ZN (N1219), .A1 (XNOR_1_3_NAND2_NUM317_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM318_OUT, XNOR_1_2_NAND2_NUM318_OUT, XNOR_1_3_NAND2_NUM318_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM318 (.ZN (XNOR_1_1_NAND2_NUM318_OUT), .A1 (N211), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM318 (.ZN (XNOR_1_2_NAND2_NUM318_OUT), .A1 (GND), .A2 (N1126));
      NOR2_X1 XNOR_1_3_NAND2_NUM318 (.ZN (XNOR_1_3_NAND2_NUM318_OUT), .A1 (XNOR_1_1_NAND2_NUM318_OUT), .A2 (XNOR_1_2_NAND2_NUM318_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM318 (.ZN (N1222), .A1 (XNOR_1_3_NAND2_NUM318_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM319_OUT, XNOR_1_2_NAND2_NUM319_OUT, XNOR_1_3_NAND2_NUM319_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM319 (.ZN (XNOR_1_1_NAND2_NUM319_OUT), .A1 (N218), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM319 (.ZN (XNOR_1_2_NAND2_NUM319_OUT), .A1 (GND), .A2 (N1129));
      NOR2_X1 XNOR_1_3_NAND2_NUM319 (.ZN (XNOR_1_3_NAND2_NUM319_OUT), .A1 (XNOR_1_1_NAND2_NUM319_OUT), .A2 (XNOR_1_2_NAND2_NUM319_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM319 (.ZN (N1225), .A1 (XNOR_1_3_NAND2_NUM319_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM320_OUT, XNOR_1_2_NAND2_NUM320_OUT, XNOR_1_3_NAND2_NUM320_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM320 (.ZN (XNOR_1_1_NAND2_NUM320_OUT), .A1 (N1), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM320 (.ZN (XNOR_1_2_NAND2_NUM320_OUT), .A1 (GND), .A2 (N1132));
      NOR2_X1 XNOR_1_3_NAND2_NUM320 (.ZN (XNOR_1_3_NAND2_NUM320_OUT), .A1 (XNOR_1_1_NAND2_NUM320_OUT), .A2 (XNOR_1_2_NAND2_NUM320_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM320 (.ZN (N1228), .A1 (XNOR_1_3_NAND2_NUM320_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM321_OUT, XNOR_1_2_NAND2_NUM321_OUT, XNOR_1_3_NAND2_NUM321_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM321 (.ZN (XNOR_1_1_NAND2_NUM321_OUT), .A1 (N1036), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM321 (.ZN (XNOR_1_2_NAND2_NUM321_OUT), .A1 (GND), .A2 (N1132));
      NOR2_X1 XNOR_1_3_NAND2_NUM321 (.ZN (XNOR_1_3_NAND2_NUM321_OUT), .A1 (XNOR_1_1_NAND2_NUM321_OUT), .A2 (XNOR_1_2_NAND2_NUM321_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM321 (.ZN (N1229), .A1 (XNOR_1_3_NAND2_NUM321_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM322_OUT, XNOR_1_2_NAND2_NUM322_OUT, XNOR_1_3_NAND2_NUM322_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM322 (.ZN (XNOR_1_1_NAND2_NUM322_OUT), .A1 (N8), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM322 (.ZN (XNOR_1_2_NAND2_NUM322_OUT), .A1 (GND), .A2 (N1135));
      NOR2_X1 XNOR_1_3_NAND2_NUM322 (.ZN (XNOR_1_3_NAND2_NUM322_OUT), .A1 (XNOR_1_1_NAND2_NUM322_OUT), .A2 (XNOR_1_2_NAND2_NUM322_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM322 (.ZN (N1230), .A1 (XNOR_1_3_NAND2_NUM322_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM323_OUT, XNOR_1_2_NAND2_NUM323_OUT, XNOR_1_3_NAND2_NUM323_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM323 (.ZN (XNOR_1_1_NAND2_NUM323_OUT), .A1 (N1039), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM323 (.ZN (XNOR_1_2_NAND2_NUM323_OUT), .A1 (GND), .A2 (N1135));
      NOR2_X1 XNOR_1_3_NAND2_NUM323 (.ZN (XNOR_1_3_NAND2_NUM323_OUT), .A1 (XNOR_1_1_NAND2_NUM323_OUT), .A2 (XNOR_1_2_NAND2_NUM323_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM323 (.ZN (N1231), .A1 (XNOR_1_3_NAND2_NUM323_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM324_OUT, XNOR_1_2_NAND2_NUM324_OUT, XNOR_1_3_NAND2_NUM324_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM324 (.ZN (XNOR_1_1_NAND2_NUM324_OUT), .A1 (N15), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM324 (.ZN (XNOR_1_2_NAND2_NUM324_OUT), .A1 (GND), .A2 (N1138));
      NOR2_X1 XNOR_1_3_NAND2_NUM324 (.ZN (XNOR_1_3_NAND2_NUM324_OUT), .A1 (XNOR_1_1_NAND2_NUM324_OUT), .A2 (XNOR_1_2_NAND2_NUM324_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM324 (.ZN (N1232), .A1 (XNOR_1_3_NAND2_NUM324_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM325_OUT, XNOR_1_2_NAND2_NUM325_OUT, XNOR_1_3_NAND2_NUM325_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM325 (.ZN (XNOR_1_1_NAND2_NUM325_OUT), .A1 (N1042), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM325 (.ZN (XNOR_1_2_NAND2_NUM325_OUT), .A1 (GND), .A2 (N1138));
      NOR2_X1 XNOR_1_3_NAND2_NUM325 (.ZN (XNOR_1_3_NAND2_NUM325_OUT), .A1 (XNOR_1_1_NAND2_NUM325_OUT), .A2 (XNOR_1_2_NAND2_NUM325_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM325 (.ZN (N1233), .A1 (XNOR_1_3_NAND2_NUM325_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM326_OUT, XNOR_1_2_NAND2_NUM326_OUT, XNOR_1_3_NAND2_NUM326_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM326 (.ZN (XNOR_1_1_NAND2_NUM326_OUT), .A1 (N22), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM326 (.ZN (XNOR_1_2_NAND2_NUM326_OUT), .A1 (GND), .A2 (N1141));
      NOR2_X1 XNOR_1_3_NAND2_NUM326 (.ZN (XNOR_1_3_NAND2_NUM326_OUT), .A1 (XNOR_1_1_NAND2_NUM326_OUT), .A2 (XNOR_1_2_NAND2_NUM326_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM326 (.ZN (N1234), .A1 (XNOR_1_3_NAND2_NUM326_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM327_OUT, XNOR_1_2_NAND2_NUM327_OUT, XNOR_1_3_NAND2_NUM327_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM327 (.ZN (XNOR_1_1_NAND2_NUM327_OUT), .A1 (N1045), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM327 (.ZN (XNOR_1_2_NAND2_NUM327_OUT), .A1 (GND), .A2 (N1141));
      NOR2_X1 XNOR_1_3_NAND2_NUM327 (.ZN (XNOR_1_3_NAND2_NUM327_OUT), .A1 (XNOR_1_1_NAND2_NUM327_OUT), .A2 (XNOR_1_2_NAND2_NUM327_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM327 (.ZN (N1235), .A1 (XNOR_1_3_NAND2_NUM327_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM328_OUT, XNOR_1_2_NAND2_NUM328_OUT, XNOR_1_3_NAND2_NUM328_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM328 (.ZN (XNOR_1_1_NAND2_NUM328_OUT), .A1 (N29), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM328 (.ZN (XNOR_1_2_NAND2_NUM328_OUT), .A1 (GND), .A2 (N1144));
      NOR2_X1 XNOR_1_3_NAND2_NUM328 (.ZN (XNOR_1_3_NAND2_NUM328_OUT), .A1 (XNOR_1_1_NAND2_NUM328_OUT), .A2 (XNOR_1_2_NAND2_NUM328_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM328 (.ZN (N1236), .A1 (XNOR_1_3_NAND2_NUM328_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM329_OUT, XNOR_1_2_NAND2_NUM329_OUT, XNOR_1_3_NAND2_NUM329_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM329 (.ZN (XNOR_1_1_NAND2_NUM329_OUT), .A1 (N1048), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM329 (.ZN (XNOR_1_2_NAND2_NUM329_OUT), .A1 (GND), .A2 (N1144));
      NOR2_X1 XNOR_1_3_NAND2_NUM329 (.ZN (XNOR_1_3_NAND2_NUM329_OUT), .A1 (XNOR_1_1_NAND2_NUM329_OUT), .A2 (XNOR_1_2_NAND2_NUM329_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM329 (.ZN (N1237), .A1 (XNOR_1_3_NAND2_NUM329_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM330_OUT, XNOR_1_2_NAND2_NUM330_OUT, XNOR_1_3_NAND2_NUM330_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM330 (.ZN (XNOR_1_1_NAND2_NUM330_OUT), .A1 (N36), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM330 (.ZN (XNOR_1_2_NAND2_NUM330_OUT), .A1 (GND), .A2 (N1147));
      NOR2_X1 XNOR_1_3_NAND2_NUM330 (.ZN (XNOR_1_3_NAND2_NUM330_OUT), .A1 (XNOR_1_1_NAND2_NUM330_OUT), .A2 (XNOR_1_2_NAND2_NUM330_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM330 (.ZN (N1238), .A1 (XNOR_1_3_NAND2_NUM330_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM331_OUT, XNOR_1_2_NAND2_NUM331_OUT, XNOR_1_3_NAND2_NUM331_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM331 (.ZN (XNOR_1_1_NAND2_NUM331_OUT), .A1 (N1051), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM331 (.ZN (XNOR_1_2_NAND2_NUM331_OUT), .A1 (GND), .A2 (N1147));
      NOR2_X1 XNOR_1_3_NAND2_NUM331 (.ZN (XNOR_1_3_NAND2_NUM331_OUT), .A1 (XNOR_1_1_NAND2_NUM331_OUT), .A2 (XNOR_1_2_NAND2_NUM331_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM331 (.ZN (N1239), .A1 (XNOR_1_3_NAND2_NUM331_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM332_OUT, XNOR_1_2_NAND2_NUM332_OUT, XNOR_1_3_NAND2_NUM332_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM332 (.ZN (XNOR_1_1_NAND2_NUM332_OUT), .A1 (N43), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM332 (.ZN (XNOR_1_2_NAND2_NUM332_OUT), .A1 (GND), .A2 (N1150));
      NOR2_X1 XNOR_1_3_NAND2_NUM332 (.ZN (XNOR_1_3_NAND2_NUM332_OUT), .A1 (XNOR_1_1_NAND2_NUM332_OUT), .A2 (XNOR_1_2_NAND2_NUM332_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM332 (.ZN (N1240), .A1 (XNOR_1_3_NAND2_NUM332_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM333_OUT, XNOR_1_2_NAND2_NUM333_OUT, XNOR_1_3_NAND2_NUM333_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM333 (.ZN (XNOR_1_1_NAND2_NUM333_OUT), .A1 (N1054), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM333 (.ZN (XNOR_1_2_NAND2_NUM333_OUT), .A1 (GND), .A2 (N1150));
      NOR2_X1 XNOR_1_3_NAND2_NUM333 (.ZN (XNOR_1_3_NAND2_NUM333_OUT), .A1 (XNOR_1_1_NAND2_NUM333_OUT), .A2 (XNOR_1_2_NAND2_NUM333_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM333 (.ZN (N1241), .A1 (XNOR_1_3_NAND2_NUM333_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM334_OUT, XNOR_1_2_NAND2_NUM334_OUT, XNOR_1_3_NAND2_NUM334_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM334 (.ZN (XNOR_1_1_NAND2_NUM334_OUT), .A1 (N50), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM334 (.ZN (XNOR_1_2_NAND2_NUM334_OUT), .A1 (GND), .A2 (N1153));
      NOR2_X1 XNOR_1_3_NAND2_NUM334 (.ZN (XNOR_1_3_NAND2_NUM334_OUT), .A1 (XNOR_1_1_NAND2_NUM334_OUT), .A2 (XNOR_1_2_NAND2_NUM334_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM334 (.ZN (N1242), .A1 (XNOR_1_3_NAND2_NUM334_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM335_OUT, XNOR_1_2_NAND2_NUM335_OUT, XNOR_1_3_NAND2_NUM335_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM335 (.ZN (XNOR_1_1_NAND2_NUM335_OUT), .A1 (N1057), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM335 (.ZN (XNOR_1_2_NAND2_NUM335_OUT), .A1 (GND), .A2 (N1153));
      NOR2_X1 XNOR_1_3_NAND2_NUM335 (.ZN (XNOR_1_3_NAND2_NUM335_OUT), .A1 (XNOR_1_1_NAND2_NUM335_OUT), .A2 (XNOR_1_2_NAND2_NUM335_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM335 (.ZN (N1243), .A1 (XNOR_1_3_NAND2_NUM335_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM336_OUT, XNOR_1_2_NAND2_NUM336_OUT, XNOR_1_3_NAND2_NUM336_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM336 (.ZN (XNOR_1_1_NAND2_NUM336_OUT), .A1 (N57), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM336 (.ZN (XNOR_1_2_NAND2_NUM336_OUT), .A1 (GND), .A2 (N1156));
      NOR2_X1 XNOR_1_3_NAND2_NUM336 (.ZN (XNOR_1_3_NAND2_NUM336_OUT), .A1 (XNOR_1_1_NAND2_NUM336_OUT), .A2 (XNOR_1_2_NAND2_NUM336_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM336 (.ZN (N1244), .A1 (XNOR_1_3_NAND2_NUM336_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM337_OUT, XNOR_1_2_NAND2_NUM337_OUT, XNOR_1_3_NAND2_NUM337_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM337 (.ZN (XNOR_1_1_NAND2_NUM337_OUT), .A1 (N1060), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM337 (.ZN (XNOR_1_2_NAND2_NUM337_OUT), .A1 (GND), .A2 (N1156));
      NOR2_X1 XNOR_1_3_NAND2_NUM337 (.ZN (XNOR_1_3_NAND2_NUM337_OUT), .A1 (XNOR_1_1_NAND2_NUM337_OUT), .A2 (XNOR_1_2_NAND2_NUM337_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM337 (.ZN (N1245), .A1 (XNOR_1_3_NAND2_NUM337_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM338_OUT, XNOR_1_2_NAND2_NUM338_OUT, XNOR_1_3_NAND2_NUM338_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM338 (.ZN (XNOR_1_1_NAND2_NUM338_OUT), .A1 (N64), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM338 (.ZN (XNOR_1_2_NAND2_NUM338_OUT), .A1 (GND), .A2 (N1159));
      NOR2_X1 XNOR_1_3_NAND2_NUM338 (.ZN (XNOR_1_3_NAND2_NUM338_OUT), .A1 (XNOR_1_1_NAND2_NUM338_OUT), .A2 (XNOR_1_2_NAND2_NUM338_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM338 (.ZN (N1246), .A1 (XNOR_1_3_NAND2_NUM338_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM339_OUT, XNOR_1_2_NAND2_NUM339_OUT, XNOR_1_3_NAND2_NUM339_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM339 (.ZN (XNOR_1_1_NAND2_NUM339_OUT), .A1 (N1063), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM339 (.ZN (XNOR_1_2_NAND2_NUM339_OUT), .A1 (GND), .A2 (N1159));
      NOR2_X1 XNOR_1_3_NAND2_NUM339 (.ZN (XNOR_1_3_NAND2_NUM339_OUT), .A1 (XNOR_1_1_NAND2_NUM339_OUT), .A2 (XNOR_1_2_NAND2_NUM339_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM339 (.ZN (N1247), .A1 (XNOR_1_3_NAND2_NUM339_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM340_OUT, XNOR_1_2_NAND2_NUM340_OUT, XNOR_1_3_NAND2_NUM340_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM340 (.ZN (XNOR_1_1_NAND2_NUM340_OUT), .A1 (N71), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM340 (.ZN (XNOR_1_2_NAND2_NUM340_OUT), .A1 (GND), .A2 (N1162));
      NOR2_X1 XNOR_1_3_NAND2_NUM340 (.ZN (XNOR_1_3_NAND2_NUM340_OUT), .A1 (XNOR_1_1_NAND2_NUM340_OUT), .A2 (XNOR_1_2_NAND2_NUM340_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM340 (.ZN (N1248), .A1 (XNOR_1_3_NAND2_NUM340_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM341_OUT, XNOR_1_2_NAND2_NUM341_OUT, XNOR_1_3_NAND2_NUM341_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM341 (.ZN (XNOR_1_1_NAND2_NUM341_OUT), .A1 (N1066), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM341 (.ZN (XNOR_1_2_NAND2_NUM341_OUT), .A1 (GND), .A2 (N1162));
      NOR2_X1 XNOR_1_3_NAND2_NUM341 (.ZN (XNOR_1_3_NAND2_NUM341_OUT), .A1 (XNOR_1_1_NAND2_NUM341_OUT), .A2 (XNOR_1_2_NAND2_NUM341_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM341 (.ZN (N1249), .A1 (XNOR_1_3_NAND2_NUM341_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM342_OUT, XNOR_1_2_NAND2_NUM342_OUT, XNOR_1_3_NAND2_NUM342_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM342 (.ZN (XNOR_1_1_NAND2_NUM342_OUT), .A1 (N78), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM342 (.ZN (XNOR_1_2_NAND2_NUM342_OUT), .A1 (GND), .A2 (N1165));
      NOR2_X1 XNOR_1_3_NAND2_NUM342 (.ZN (XNOR_1_3_NAND2_NUM342_OUT), .A1 (XNOR_1_1_NAND2_NUM342_OUT), .A2 (XNOR_1_2_NAND2_NUM342_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM342 (.ZN (N1250), .A1 (XNOR_1_3_NAND2_NUM342_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM343_OUT, XNOR_1_2_NAND2_NUM343_OUT, XNOR_1_3_NAND2_NUM343_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM343 (.ZN (XNOR_1_1_NAND2_NUM343_OUT), .A1 (N1069), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM343 (.ZN (XNOR_1_2_NAND2_NUM343_OUT), .A1 (GND), .A2 (N1165));
      NOR2_X1 XNOR_1_3_NAND2_NUM343 (.ZN (XNOR_1_3_NAND2_NUM343_OUT), .A1 (XNOR_1_1_NAND2_NUM343_OUT), .A2 (XNOR_1_2_NAND2_NUM343_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM343 (.ZN (N1251), .A1 (XNOR_1_3_NAND2_NUM343_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM344_OUT, XNOR_1_2_NAND2_NUM344_OUT, XNOR_1_3_NAND2_NUM344_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM344 (.ZN (XNOR_1_1_NAND2_NUM344_OUT), .A1 (N85), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM344 (.ZN (XNOR_1_2_NAND2_NUM344_OUT), .A1 (GND), .A2 (N1168));
      NOR2_X1 XNOR_1_3_NAND2_NUM344 (.ZN (XNOR_1_3_NAND2_NUM344_OUT), .A1 (XNOR_1_1_NAND2_NUM344_OUT), .A2 (XNOR_1_2_NAND2_NUM344_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM344 (.ZN (N1252), .A1 (XNOR_1_3_NAND2_NUM344_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM345_OUT, XNOR_1_2_NAND2_NUM345_OUT, XNOR_1_3_NAND2_NUM345_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM345 (.ZN (XNOR_1_1_NAND2_NUM345_OUT), .A1 (N1072), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM345 (.ZN (XNOR_1_2_NAND2_NUM345_OUT), .A1 (GND), .A2 (N1168));
      NOR2_X1 XNOR_1_3_NAND2_NUM345 (.ZN (XNOR_1_3_NAND2_NUM345_OUT), .A1 (XNOR_1_1_NAND2_NUM345_OUT), .A2 (XNOR_1_2_NAND2_NUM345_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM345 (.ZN (N1253), .A1 (XNOR_1_3_NAND2_NUM345_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM346_OUT, XNOR_1_2_NAND2_NUM346_OUT, XNOR_1_3_NAND2_NUM346_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM346 (.ZN (XNOR_1_1_NAND2_NUM346_OUT), .A1 (N92), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM346 (.ZN (XNOR_1_2_NAND2_NUM346_OUT), .A1 (GND), .A2 (N1171));
      NOR2_X1 XNOR_1_3_NAND2_NUM346 (.ZN (XNOR_1_3_NAND2_NUM346_OUT), .A1 (XNOR_1_1_NAND2_NUM346_OUT), .A2 (XNOR_1_2_NAND2_NUM346_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM346 (.ZN (N1254), .A1 (XNOR_1_3_NAND2_NUM346_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM347_OUT, XNOR_1_2_NAND2_NUM347_OUT, XNOR_1_3_NAND2_NUM347_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM347 (.ZN (XNOR_1_1_NAND2_NUM347_OUT), .A1 (N1075), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM347 (.ZN (XNOR_1_2_NAND2_NUM347_OUT), .A1 (GND), .A2 (N1171));
      NOR2_X1 XNOR_1_3_NAND2_NUM347 (.ZN (XNOR_1_3_NAND2_NUM347_OUT), .A1 (XNOR_1_1_NAND2_NUM347_OUT), .A2 (XNOR_1_2_NAND2_NUM347_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM347 (.ZN (N1255), .A1 (XNOR_1_3_NAND2_NUM347_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM348_OUT, XNOR_1_2_NAND2_NUM348_OUT, XNOR_1_3_NAND2_NUM348_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM348 (.ZN (XNOR_1_1_NAND2_NUM348_OUT), .A1 (N99), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM348 (.ZN (XNOR_1_2_NAND2_NUM348_OUT), .A1 (GND), .A2 (N1174));
      NOR2_X1 XNOR_1_3_NAND2_NUM348 (.ZN (XNOR_1_3_NAND2_NUM348_OUT), .A1 (XNOR_1_1_NAND2_NUM348_OUT), .A2 (XNOR_1_2_NAND2_NUM348_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM348 (.ZN (N1256), .A1 (XNOR_1_3_NAND2_NUM348_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM349_OUT, XNOR_1_2_NAND2_NUM349_OUT, XNOR_1_3_NAND2_NUM349_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM349 (.ZN (XNOR_1_1_NAND2_NUM349_OUT), .A1 (N1078), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM349 (.ZN (XNOR_1_2_NAND2_NUM349_OUT), .A1 (GND), .A2 (N1174));
      NOR2_X1 XNOR_1_3_NAND2_NUM349 (.ZN (XNOR_1_3_NAND2_NUM349_OUT), .A1 (XNOR_1_1_NAND2_NUM349_OUT), .A2 (XNOR_1_2_NAND2_NUM349_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM349 (.ZN (N1257), .A1 (XNOR_1_3_NAND2_NUM349_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM350_OUT, XNOR_1_2_NAND2_NUM350_OUT, XNOR_1_3_NAND2_NUM350_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM350 (.ZN (XNOR_1_1_NAND2_NUM350_OUT), .A1 (N106), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM350 (.ZN (XNOR_1_2_NAND2_NUM350_OUT), .A1 (GND), .A2 (N1177));
      NOR2_X1 XNOR_1_3_NAND2_NUM350 (.ZN (XNOR_1_3_NAND2_NUM350_OUT), .A1 (XNOR_1_1_NAND2_NUM350_OUT), .A2 (XNOR_1_2_NAND2_NUM350_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM350 (.ZN (N1258), .A1 (XNOR_1_3_NAND2_NUM350_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM351_OUT, XNOR_1_2_NAND2_NUM351_OUT, XNOR_1_3_NAND2_NUM351_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM351 (.ZN (XNOR_1_1_NAND2_NUM351_OUT), .A1 (N1081), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM351 (.ZN (XNOR_1_2_NAND2_NUM351_OUT), .A1 (GND), .A2 (N1177));
      NOR2_X1 XNOR_1_3_NAND2_NUM351 (.ZN (XNOR_1_3_NAND2_NUM351_OUT), .A1 (XNOR_1_1_NAND2_NUM351_OUT), .A2 (XNOR_1_2_NAND2_NUM351_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM351 (.ZN (N1259), .A1 (XNOR_1_3_NAND2_NUM351_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM352_OUT, XNOR_1_2_NAND2_NUM352_OUT, XNOR_1_3_NAND2_NUM352_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM352 (.ZN (XNOR_1_1_NAND2_NUM352_OUT), .A1 (N113), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM352 (.ZN (XNOR_1_2_NAND2_NUM352_OUT), .A1 (GND), .A2 (N1180));
      NOR2_X1 XNOR_1_3_NAND2_NUM352 (.ZN (XNOR_1_3_NAND2_NUM352_OUT), .A1 (XNOR_1_1_NAND2_NUM352_OUT), .A2 (XNOR_1_2_NAND2_NUM352_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM352 (.ZN (N1260), .A1 (XNOR_1_3_NAND2_NUM352_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM353_OUT, XNOR_1_2_NAND2_NUM353_OUT, XNOR_1_3_NAND2_NUM353_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM353 (.ZN (XNOR_1_1_NAND2_NUM353_OUT), .A1 (N1084), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM353 (.ZN (XNOR_1_2_NAND2_NUM353_OUT), .A1 (GND), .A2 (N1180));
      NOR2_X1 XNOR_1_3_NAND2_NUM353 (.ZN (XNOR_1_3_NAND2_NUM353_OUT), .A1 (XNOR_1_1_NAND2_NUM353_OUT), .A2 (XNOR_1_2_NAND2_NUM353_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM353 (.ZN (N1261), .A1 (XNOR_1_3_NAND2_NUM353_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM354_OUT, XNOR_1_2_NAND2_NUM354_OUT, XNOR_1_3_NAND2_NUM354_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM354 (.ZN (XNOR_1_1_NAND2_NUM354_OUT), .A1 (N120), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM354 (.ZN (XNOR_1_2_NAND2_NUM354_OUT), .A1 (GND), .A2 (N1183));
      NOR2_X1 XNOR_1_3_NAND2_NUM354 (.ZN (XNOR_1_3_NAND2_NUM354_OUT), .A1 (XNOR_1_1_NAND2_NUM354_OUT), .A2 (XNOR_1_2_NAND2_NUM354_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM354 (.ZN (N1262), .A1 (XNOR_1_3_NAND2_NUM354_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM355_OUT, XNOR_1_2_NAND2_NUM355_OUT, XNOR_1_3_NAND2_NUM355_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM355 (.ZN (XNOR_1_1_NAND2_NUM355_OUT), .A1 (N1087), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM355 (.ZN (XNOR_1_2_NAND2_NUM355_OUT), .A1 (GND), .A2 (N1183));
      NOR2_X1 XNOR_1_3_NAND2_NUM355 (.ZN (XNOR_1_3_NAND2_NUM355_OUT), .A1 (XNOR_1_1_NAND2_NUM355_OUT), .A2 (XNOR_1_2_NAND2_NUM355_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM355 (.ZN (N1263), .A1 (XNOR_1_3_NAND2_NUM355_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM356_OUT, XNOR_1_2_NAND2_NUM356_OUT, XNOR_1_3_NAND2_NUM356_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM356 (.ZN (XNOR_1_1_NAND2_NUM356_OUT), .A1 (N127), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM356 (.ZN (XNOR_1_2_NAND2_NUM356_OUT), .A1 (GND), .A2 (N1186));
      NOR2_X1 XNOR_1_3_NAND2_NUM356 (.ZN (XNOR_1_3_NAND2_NUM356_OUT), .A1 (XNOR_1_1_NAND2_NUM356_OUT), .A2 (XNOR_1_2_NAND2_NUM356_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM356 (.ZN (N1264), .A1 (XNOR_1_3_NAND2_NUM356_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM357_OUT, XNOR_1_2_NAND2_NUM357_OUT, XNOR_1_3_NAND2_NUM357_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM357 (.ZN (XNOR_1_1_NAND2_NUM357_OUT), .A1 (N1090), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM357 (.ZN (XNOR_1_2_NAND2_NUM357_OUT), .A1 (GND), .A2 (N1186));
      NOR2_X1 XNOR_1_3_NAND2_NUM357 (.ZN (XNOR_1_3_NAND2_NUM357_OUT), .A1 (XNOR_1_1_NAND2_NUM357_OUT), .A2 (XNOR_1_2_NAND2_NUM357_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM357 (.ZN (N1265), .A1 (XNOR_1_3_NAND2_NUM357_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM358_OUT, XNOR_1_2_NAND2_NUM358_OUT, XNOR_1_3_NAND2_NUM358_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM358 (.ZN (XNOR_1_1_NAND2_NUM358_OUT), .A1 (N134), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM358 (.ZN (XNOR_1_2_NAND2_NUM358_OUT), .A1 (GND), .A2 (N1189));
      NOR2_X1 XNOR_1_3_NAND2_NUM358 (.ZN (XNOR_1_3_NAND2_NUM358_OUT), .A1 (XNOR_1_1_NAND2_NUM358_OUT), .A2 (XNOR_1_2_NAND2_NUM358_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM358 (.ZN (N1266), .A1 (XNOR_1_3_NAND2_NUM358_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM359_OUT, XNOR_1_2_NAND2_NUM359_OUT, XNOR_1_3_NAND2_NUM359_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM359 (.ZN (XNOR_1_1_NAND2_NUM359_OUT), .A1 (N1093), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM359 (.ZN (XNOR_1_2_NAND2_NUM359_OUT), .A1 (GND), .A2 (N1189));
      NOR2_X1 XNOR_1_3_NAND2_NUM359 (.ZN (XNOR_1_3_NAND2_NUM359_OUT), .A1 (XNOR_1_1_NAND2_NUM359_OUT), .A2 (XNOR_1_2_NAND2_NUM359_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM359 (.ZN (N1267), .A1 (XNOR_1_3_NAND2_NUM359_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM360_OUT, XNOR_1_2_NAND2_NUM360_OUT, XNOR_1_3_NAND2_NUM360_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM360 (.ZN (XNOR_1_1_NAND2_NUM360_OUT), .A1 (N141), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM360 (.ZN (XNOR_1_2_NAND2_NUM360_OUT), .A1 (GND), .A2 (N1192));
      NOR2_X1 XNOR_1_3_NAND2_NUM360 (.ZN (XNOR_1_3_NAND2_NUM360_OUT), .A1 (XNOR_1_1_NAND2_NUM360_OUT), .A2 (XNOR_1_2_NAND2_NUM360_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM360 (.ZN (N1268), .A1 (XNOR_1_3_NAND2_NUM360_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM361_OUT, XNOR_1_2_NAND2_NUM361_OUT, XNOR_1_3_NAND2_NUM361_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM361 (.ZN (XNOR_1_1_NAND2_NUM361_OUT), .A1 (N1096), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM361 (.ZN (XNOR_1_2_NAND2_NUM361_OUT), .A1 (GND), .A2 (N1192));
      NOR2_X1 XNOR_1_3_NAND2_NUM361 (.ZN (XNOR_1_3_NAND2_NUM361_OUT), .A1 (XNOR_1_1_NAND2_NUM361_OUT), .A2 (XNOR_1_2_NAND2_NUM361_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM361 (.ZN (N1269), .A1 (XNOR_1_3_NAND2_NUM361_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM362_OUT, XNOR_1_2_NAND2_NUM362_OUT, XNOR_1_3_NAND2_NUM362_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM362 (.ZN (XNOR_1_1_NAND2_NUM362_OUT), .A1 (N148), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM362 (.ZN (XNOR_1_2_NAND2_NUM362_OUT), .A1 (GND), .A2 (N1195));
      NOR2_X1 XNOR_1_3_NAND2_NUM362 (.ZN (XNOR_1_3_NAND2_NUM362_OUT), .A1 (XNOR_1_1_NAND2_NUM362_OUT), .A2 (XNOR_1_2_NAND2_NUM362_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM362 (.ZN (N1270), .A1 (XNOR_1_3_NAND2_NUM362_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM363_OUT, XNOR_1_2_NAND2_NUM363_OUT, XNOR_1_3_NAND2_NUM363_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM363 (.ZN (XNOR_1_1_NAND2_NUM363_OUT), .A1 (N1099), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM363 (.ZN (XNOR_1_2_NAND2_NUM363_OUT), .A1 (GND), .A2 (N1195));
      NOR2_X1 XNOR_1_3_NAND2_NUM363 (.ZN (XNOR_1_3_NAND2_NUM363_OUT), .A1 (XNOR_1_1_NAND2_NUM363_OUT), .A2 (XNOR_1_2_NAND2_NUM363_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM363 (.ZN (N1271), .A1 (XNOR_1_3_NAND2_NUM363_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM364_OUT, XNOR_1_2_NAND2_NUM364_OUT, XNOR_1_3_NAND2_NUM364_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM364 (.ZN (XNOR_1_1_NAND2_NUM364_OUT), .A1 (N155), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM364 (.ZN (XNOR_1_2_NAND2_NUM364_OUT), .A1 (GND), .A2 (N1198));
      NOR2_X1 XNOR_1_3_NAND2_NUM364 (.ZN (XNOR_1_3_NAND2_NUM364_OUT), .A1 (XNOR_1_1_NAND2_NUM364_OUT), .A2 (XNOR_1_2_NAND2_NUM364_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM364 (.ZN (N1272), .A1 (XNOR_1_3_NAND2_NUM364_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM365_OUT, XNOR_1_2_NAND2_NUM365_OUT, XNOR_1_3_NAND2_NUM365_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM365 (.ZN (XNOR_1_1_NAND2_NUM365_OUT), .A1 (N1102), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM365 (.ZN (XNOR_1_2_NAND2_NUM365_OUT), .A1 (GND), .A2 (N1198));
      NOR2_X1 XNOR_1_3_NAND2_NUM365 (.ZN (XNOR_1_3_NAND2_NUM365_OUT), .A1 (XNOR_1_1_NAND2_NUM365_OUT), .A2 (XNOR_1_2_NAND2_NUM365_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM365 (.ZN (N1273), .A1 (XNOR_1_3_NAND2_NUM365_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM366_OUT, XNOR_1_2_NAND2_NUM366_OUT, XNOR_1_3_NAND2_NUM366_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM366 (.ZN (XNOR_1_1_NAND2_NUM366_OUT), .A1 (N162), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM366 (.ZN (XNOR_1_2_NAND2_NUM366_OUT), .A1 (GND), .A2 (N1201));
      NOR2_X1 XNOR_1_3_NAND2_NUM366 (.ZN (XNOR_1_3_NAND2_NUM366_OUT), .A1 (XNOR_1_1_NAND2_NUM366_OUT), .A2 (XNOR_1_2_NAND2_NUM366_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM366 (.ZN (N1274), .A1 (XNOR_1_3_NAND2_NUM366_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM367_OUT, XNOR_1_2_NAND2_NUM367_OUT, XNOR_1_3_NAND2_NUM367_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM367 (.ZN (XNOR_1_1_NAND2_NUM367_OUT), .A1 (N1105), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM367 (.ZN (XNOR_1_2_NAND2_NUM367_OUT), .A1 (GND), .A2 (N1201));
      NOR2_X1 XNOR_1_3_NAND2_NUM367 (.ZN (XNOR_1_3_NAND2_NUM367_OUT), .A1 (XNOR_1_1_NAND2_NUM367_OUT), .A2 (XNOR_1_2_NAND2_NUM367_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM367 (.ZN (N1275), .A1 (XNOR_1_3_NAND2_NUM367_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM368_OUT, XNOR_1_2_NAND2_NUM368_OUT, XNOR_1_3_NAND2_NUM368_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM368 (.ZN (XNOR_1_1_NAND2_NUM368_OUT), .A1 (N169), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM368 (.ZN (XNOR_1_2_NAND2_NUM368_OUT), .A1 (GND), .A2 (N1204));
      NOR2_X1 XNOR_1_3_NAND2_NUM368 (.ZN (XNOR_1_3_NAND2_NUM368_OUT), .A1 (XNOR_1_1_NAND2_NUM368_OUT), .A2 (XNOR_1_2_NAND2_NUM368_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM368 (.ZN (N1276), .A1 (XNOR_1_3_NAND2_NUM368_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM369_OUT, XNOR_1_2_NAND2_NUM369_OUT, XNOR_1_3_NAND2_NUM369_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM369 (.ZN (XNOR_1_1_NAND2_NUM369_OUT), .A1 (N1108), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM369 (.ZN (XNOR_1_2_NAND2_NUM369_OUT), .A1 (GND), .A2 (N1204));
      NOR2_X1 XNOR_1_3_NAND2_NUM369 (.ZN (XNOR_1_3_NAND2_NUM369_OUT), .A1 (XNOR_1_1_NAND2_NUM369_OUT), .A2 (XNOR_1_2_NAND2_NUM369_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM369 (.ZN (N1277), .A1 (XNOR_1_3_NAND2_NUM369_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM370_OUT, XNOR_1_2_NAND2_NUM370_OUT, XNOR_1_3_NAND2_NUM370_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM370 (.ZN (XNOR_1_1_NAND2_NUM370_OUT), .A1 (N176), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM370 (.ZN (XNOR_1_2_NAND2_NUM370_OUT), .A1 (GND), .A2 (N1207));
      NOR2_X1 XNOR_1_3_NAND2_NUM370 (.ZN (XNOR_1_3_NAND2_NUM370_OUT), .A1 (XNOR_1_1_NAND2_NUM370_OUT), .A2 (XNOR_1_2_NAND2_NUM370_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM370 (.ZN (N1278), .A1 (XNOR_1_3_NAND2_NUM370_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM371_OUT, XNOR_1_2_NAND2_NUM371_OUT, XNOR_1_3_NAND2_NUM371_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM371 (.ZN (XNOR_1_1_NAND2_NUM371_OUT), .A1 (N1111), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM371 (.ZN (XNOR_1_2_NAND2_NUM371_OUT), .A1 (GND), .A2 (N1207));
      NOR2_X1 XNOR_1_3_NAND2_NUM371 (.ZN (XNOR_1_3_NAND2_NUM371_OUT), .A1 (XNOR_1_1_NAND2_NUM371_OUT), .A2 (XNOR_1_2_NAND2_NUM371_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM371 (.ZN (N1279), .A1 (XNOR_1_3_NAND2_NUM371_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM372_OUT, XNOR_1_2_NAND2_NUM372_OUT, XNOR_1_3_NAND2_NUM372_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM372 (.ZN (XNOR_1_1_NAND2_NUM372_OUT), .A1 (N183), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM372 (.ZN (XNOR_1_2_NAND2_NUM372_OUT), .A1 (GND), .A2 (N1210));
      NOR2_X1 XNOR_1_3_NAND2_NUM372 (.ZN (XNOR_1_3_NAND2_NUM372_OUT), .A1 (XNOR_1_1_NAND2_NUM372_OUT), .A2 (XNOR_1_2_NAND2_NUM372_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM372 (.ZN (N1280), .A1 (XNOR_1_3_NAND2_NUM372_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM373_OUT, XNOR_1_2_NAND2_NUM373_OUT, XNOR_1_3_NAND2_NUM373_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM373 (.ZN (XNOR_1_1_NAND2_NUM373_OUT), .A1 (N1114), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM373 (.ZN (XNOR_1_2_NAND2_NUM373_OUT), .A1 (GND), .A2 (N1210));
      NOR2_X1 XNOR_1_3_NAND2_NUM373 (.ZN (XNOR_1_3_NAND2_NUM373_OUT), .A1 (XNOR_1_1_NAND2_NUM373_OUT), .A2 (XNOR_1_2_NAND2_NUM373_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM373 (.ZN (N1281), .A1 (XNOR_1_3_NAND2_NUM373_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM374_OUT, XNOR_1_2_NAND2_NUM374_OUT, XNOR_1_3_NAND2_NUM374_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM374 (.ZN (XNOR_1_1_NAND2_NUM374_OUT), .A1 (N190), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM374 (.ZN (XNOR_1_2_NAND2_NUM374_OUT), .A1 (GND), .A2 (N1213));
      NOR2_X1 XNOR_1_3_NAND2_NUM374 (.ZN (XNOR_1_3_NAND2_NUM374_OUT), .A1 (XNOR_1_1_NAND2_NUM374_OUT), .A2 (XNOR_1_2_NAND2_NUM374_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM374 (.ZN (N1282), .A1 (XNOR_1_3_NAND2_NUM374_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM375_OUT, XNOR_1_2_NAND2_NUM375_OUT, XNOR_1_3_NAND2_NUM375_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM375 (.ZN (XNOR_1_1_NAND2_NUM375_OUT), .A1 (N1117), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM375 (.ZN (XNOR_1_2_NAND2_NUM375_OUT), .A1 (GND), .A2 (N1213));
      NOR2_X1 XNOR_1_3_NAND2_NUM375 (.ZN (XNOR_1_3_NAND2_NUM375_OUT), .A1 (XNOR_1_1_NAND2_NUM375_OUT), .A2 (XNOR_1_2_NAND2_NUM375_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM375 (.ZN (N1283), .A1 (XNOR_1_3_NAND2_NUM375_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM376_OUT, XNOR_1_2_NAND2_NUM376_OUT, XNOR_1_3_NAND2_NUM376_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM376 (.ZN (XNOR_1_1_NAND2_NUM376_OUT), .A1 (N197), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM376 (.ZN (XNOR_1_2_NAND2_NUM376_OUT), .A1 (GND), .A2 (N1216));
      NOR2_X1 XNOR_1_3_NAND2_NUM376 (.ZN (XNOR_1_3_NAND2_NUM376_OUT), .A1 (XNOR_1_1_NAND2_NUM376_OUT), .A2 (XNOR_1_2_NAND2_NUM376_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM376 (.ZN (N1284), .A1 (XNOR_1_3_NAND2_NUM376_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM377_OUT, XNOR_1_2_NAND2_NUM377_OUT, XNOR_1_3_NAND2_NUM377_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM377 (.ZN (XNOR_1_1_NAND2_NUM377_OUT), .A1 (N1120), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM377 (.ZN (XNOR_1_2_NAND2_NUM377_OUT), .A1 (GND), .A2 (N1216));
      NOR2_X1 XNOR_1_3_NAND2_NUM377 (.ZN (XNOR_1_3_NAND2_NUM377_OUT), .A1 (XNOR_1_1_NAND2_NUM377_OUT), .A2 (XNOR_1_2_NAND2_NUM377_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM377 (.ZN (N1285), .A1 (XNOR_1_3_NAND2_NUM377_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM378_OUT, XNOR_1_2_NAND2_NUM378_OUT, XNOR_1_3_NAND2_NUM378_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM378 (.ZN (XNOR_1_1_NAND2_NUM378_OUT), .A1 (N204), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM378 (.ZN (XNOR_1_2_NAND2_NUM378_OUT), .A1 (GND), .A2 (N1219));
      NOR2_X1 XNOR_1_3_NAND2_NUM378 (.ZN (XNOR_1_3_NAND2_NUM378_OUT), .A1 (XNOR_1_1_NAND2_NUM378_OUT), .A2 (XNOR_1_2_NAND2_NUM378_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM378 (.ZN (N1286), .A1 (XNOR_1_3_NAND2_NUM378_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM379_OUT, XNOR_1_2_NAND2_NUM379_OUT, XNOR_1_3_NAND2_NUM379_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM379 (.ZN (XNOR_1_1_NAND2_NUM379_OUT), .A1 (N1123), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM379 (.ZN (XNOR_1_2_NAND2_NUM379_OUT), .A1 (GND), .A2 (N1219));
      NOR2_X1 XNOR_1_3_NAND2_NUM379 (.ZN (XNOR_1_3_NAND2_NUM379_OUT), .A1 (XNOR_1_1_NAND2_NUM379_OUT), .A2 (XNOR_1_2_NAND2_NUM379_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM379 (.ZN (N1287), .A1 (XNOR_1_3_NAND2_NUM379_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM380_OUT, XNOR_1_2_NAND2_NUM380_OUT, XNOR_1_3_NAND2_NUM380_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM380 (.ZN (XNOR_1_1_NAND2_NUM380_OUT), .A1 (N211), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM380 (.ZN (XNOR_1_2_NAND2_NUM380_OUT), .A1 (GND), .A2 (N1222));
      NOR2_X1 XNOR_1_3_NAND2_NUM380 (.ZN (XNOR_1_3_NAND2_NUM380_OUT), .A1 (XNOR_1_1_NAND2_NUM380_OUT), .A2 (XNOR_1_2_NAND2_NUM380_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM380 (.ZN (N1288), .A1 (XNOR_1_3_NAND2_NUM380_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM381_OUT, XNOR_1_2_NAND2_NUM381_OUT, XNOR_1_3_NAND2_NUM381_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM381 (.ZN (XNOR_1_1_NAND2_NUM381_OUT), .A1 (N1126), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM381 (.ZN (XNOR_1_2_NAND2_NUM381_OUT), .A1 (GND), .A2 (N1222));
      NOR2_X1 XNOR_1_3_NAND2_NUM381 (.ZN (XNOR_1_3_NAND2_NUM381_OUT), .A1 (XNOR_1_1_NAND2_NUM381_OUT), .A2 (XNOR_1_2_NAND2_NUM381_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM381 (.ZN (N1289), .A1 (XNOR_1_3_NAND2_NUM381_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM382_OUT, XNOR_1_2_NAND2_NUM382_OUT, XNOR_1_3_NAND2_NUM382_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM382 (.ZN (XNOR_1_1_NAND2_NUM382_OUT), .A1 (N218), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM382 (.ZN (XNOR_1_2_NAND2_NUM382_OUT), .A1 (GND), .A2 (N1225));
      NOR2_X1 XNOR_1_3_NAND2_NUM382 (.ZN (XNOR_1_3_NAND2_NUM382_OUT), .A1 (XNOR_1_1_NAND2_NUM382_OUT), .A2 (XNOR_1_2_NAND2_NUM382_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM382 (.ZN (N1290), .A1 (XNOR_1_3_NAND2_NUM382_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM383_OUT, XNOR_1_2_NAND2_NUM383_OUT, XNOR_1_3_NAND2_NUM383_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM383 (.ZN (XNOR_1_1_NAND2_NUM383_OUT), .A1 (N1129), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM383 (.ZN (XNOR_1_2_NAND2_NUM383_OUT), .A1 (GND), .A2 (N1225));
      NOR2_X1 XNOR_1_3_NAND2_NUM383 (.ZN (XNOR_1_3_NAND2_NUM383_OUT), .A1 (XNOR_1_1_NAND2_NUM383_OUT), .A2 (XNOR_1_2_NAND2_NUM383_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM383 (.ZN (N1291), .A1 (XNOR_1_3_NAND2_NUM383_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM384_OUT, XNOR_1_2_NAND2_NUM384_OUT, XNOR_1_3_NAND2_NUM384_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM384 (.ZN (XNOR_1_1_NAND2_NUM384_OUT), .A1 (N1228), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM384 (.ZN (XNOR_1_2_NAND2_NUM384_OUT), .A1 (GND), .A2 (N1229));
      NOR2_X1 XNOR_1_3_NAND2_NUM384 (.ZN (XNOR_1_3_NAND2_NUM384_OUT), .A1 (XNOR_1_1_NAND2_NUM384_OUT), .A2 (XNOR_1_2_NAND2_NUM384_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM384 (.ZN (N1292), .A1 (XNOR_1_3_NAND2_NUM384_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM385_OUT, XNOR_1_2_NAND2_NUM385_OUT, XNOR_1_3_NAND2_NUM385_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM385 (.ZN (XNOR_1_1_NAND2_NUM385_OUT), .A1 (N1230), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM385 (.ZN (XNOR_1_2_NAND2_NUM385_OUT), .A1 (GND), .A2 (N1231));
      NOR2_X1 XNOR_1_3_NAND2_NUM385 (.ZN (XNOR_1_3_NAND2_NUM385_OUT), .A1 (XNOR_1_1_NAND2_NUM385_OUT), .A2 (XNOR_1_2_NAND2_NUM385_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM385 (.ZN (N1293), .A1 (XNOR_1_3_NAND2_NUM385_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM386_OUT, XNOR_1_2_NAND2_NUM386_OUT, XNOR_1_3_NAND2_NUM386_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM386 (.ZN (XNOR_1_1_NAND2_NUM386_OUT), .A1 (N1232), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM386 (.ZN (XNOR_1_2_NAND2_NUM386_OUT), .A1 (GND), .A2 (N1233));
      NOR2_X1 XNOR_1_3_NAND2_NUM386 (.ZN (XNOR_1_3_NAND2_NUM386_OUT), .A1 (XNOR_1_1_NAND2_NUM386_OUT), .A2 (XNOR_1_2_NAND2_NUM386_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM386 (.ZN (N1294), .A1 (XNOR_1_3_NAND2_NUM386_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM387_OUT, XNOR_1_2_NAND2_NUM387_OUT, XNOR_1_3_NAND2_NUM387_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM387 (.ZN (XNOR_1_1_NAND2_NUM387_OUT), .A1 (N1234), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM387 (.ZN (XNOR_1_2_NAND2_NUM387_OUT), .A1 (GND), .A2 (N1235));
      NOR2_X1 XNOR_1_3_NAND2_NUM387 (.ZN (XNOR_1_3_NAND2_NUM387_OUT), .A1 (XNOR_1_1_NAND2_NUM387_OUT), .A2 (XNOR_1_2_NAND2_NUM387_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM387 (.ZN (N1295), .A1 (XNOR_1_3_NAND2_NUM387_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM388_OUT, XNOR_1_2_NAND2_NUM388_OUT, XNOR_1_3_NAND2_NUM388_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM388 (.ZN (XNOR_1_1_NAND2_NUM388_OUT), .A1 (N1236), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM388 (.ZN (XNOR_1_2_NAND2_NUM388_OUT), .A1 (GND), .A2 (N1237));
      NOR2_X1 XNOR_1_3_NAND2_NUM388 (.ZN (XNOR_1_3_NAND2_NUM388_OUT), .A1 (XNOR_1_1_NAND2_NUM388_OUT), .A2 (XNOR_1_2_NAND2_NUM388_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM388 (.ZN (N1296), .A1 (XNOR_1_3_NAND2_NUM388_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM389_OUT, XNOR_1_2_NAND2_NUM389_OUT, XNOR_1_3_NAND2_NUM389_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM389 (.ZN (XNOR_1_1_NAND2_NUM389_OUT), .A1 (N1238), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM389 (.ZN (XNOR_1_2_NAND2_NUM389_OUT), .A1 (GND), .A2 (N1239));
      NOR2_X1 XNOR_1_3_NAND2_NUM389 (.ZN (XNOR_1_3_NAND2_NUM389_OUT), .A1 (XNOR_1_1_NAND2_NUM389_OUT), .A2 (XNOR_1_2_NAND2_NUM389_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM389 (.ZN (N1297), .A1 (XNOR_1_3_NAND2_NUM389_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM390_OUT, XNOR_1_2_NAND2_NUM390_OUT, XNOR_1_3_NAND2_NUM390_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM390 (.ZN (XNOR_1_1_NAND2_NUM390_OUT), .A1 (N1240), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM390 (.ZN (XNOR_1_2_NAND2_NUM390_OUT), .A1 (GND), .A2 (N1241));
      NOR2_X1 XNOR_1_3_NAND2_NUM390 (.ZN (XNOR_1_3_NAND2_NUM390_OUT), .A1 (XNOR_1_1_NAND2_NUM390_OUT), .A2 (XNOR_1_2_NAND2_NUM390_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM390 (.ZN (N1298), .A1 (XNOR_1_3_NAND2_NUM390_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM391_OUT, XNOR_1_2_NAND2_NUM391_OUT, XNOR_1_3_NAND2_NUM391_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM391 (.ZN (XNOR_1_1_NAND2_NUM391_OUT), .A1 (N1242), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM391 (.ZN (XNOR_1_2_NAND2_NUM391_OUT), .A1 (GND), .A2 (N1243));
      NOR2_X1 XNOR_1_3_NAND2_NUM391 (.ZN (XNOR_1_3_NAND2_NUM391_OUT), .A1 (XNOR_1_1_NAND2_NUM391_OUT), .A2 (XNOR_1_2_NAND2_NUM391_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM391 (.ZN (N1299), .A1 (XNOR_1_3_NAND2_NUM391_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM392_OUT, XNOR_1_2_NAND2_NUM392_OUT, XNOR_1_3_NAND2_NUM392_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM392 (.ZN (XNOR_1_1_NAND2_NUM392_OUT), .A1 (N1244), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM392 (.ZN (XNOR_1_2_NAND2_NUM392_OUT), .A1 (GND), .A2 (N1245));
      NOR2_X1 XNOR_1_3_NAND2_NUM392 (.ZN (XNOR_1_3_NAND2_NUM392_OUT), .A1 (XNOR_1_1_NAND2_NUM392_OUT), .A2 (XNOR_1_2_NAND2_NUM392_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM392 (.ZN (N1300), .A1 (XNOR_1_3_NAND2_NUM392_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM393_OUT, XNOR_1_2_NAND2_NUM393_OUT, XNOR_1_3_NAND2_NUM393_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM393 (.ZN (XNOR_1_1_NAND2_NUM393_OUT), .A1 (N1246), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM393 (.ZN (XNOR_1_2_NAND2_NUM393_OUT), .A1 (GND), .A2 (N1247));
      NOR2_X1 XNOR_1_3_NAND2_NUM393 (.ZN (XNOR_1_3_NAND2_NUM393_OUT), .A1 (XNOR_1_1_NAND2_NUM393_OUT), .A2 (XNOR_1_2_NAND2_NUM393_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM393 (.ZN (N1301), .A1 (XNOR_1_3_NAND2_NUM393_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM394_OUT, XNOR_1_2_NAND2_NUM394_OUT, XNOR_1_3_NAND2_NUM394_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM394 (.ZN (XNOR_1_1_NAND2_NUM394_OUT), .A1 (N1248), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM394 (.ZN (XNOR_1_2_NAND2_NUM394_OUT), .A1 (GND), .A2 (N1249));
      NOR2_X1 XNOR_1_3_NAND2_NUM394 (.ZN (XNOR_1_3_NAND2_NUM394_OUT), .A1 (XNOR_1_1_NAND2_NUM394_OUT), .A2 (XNOR_1_2_NAND2_NUM394_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM394 (.ZN (N1302), .A1 (XNOR_1_3_NAND2_NUM394_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM395_OUT, XNOR_1_2_NAND2_NUM395_OUT, XNOR_1_3_NAND2_NUM395_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM395 (.ZN (XNOR_1_1_NAND2_NUM395_OUT), .A1 (N1250), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM395 (.ZN (XNOR_1_2_NAND2_NUM395_OUT), .A1 (GND), .A2 (N1251));
      NOR2_X1 XNOR_1_3_NAND2_NUM395 (.ZN (XNOR_1_3_NAND2_NUM395_OUT), .A1 (XNOR_1_1_NAND2_NUM395_OUT), .A2 (XNOR_1_2_NAND2_NUM395_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM395 (.ZN (N1303), .A1 (XNOR_1_3_NAND2_NUM395_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM396_OUT, XNOR_1_2_NAND2_NUM396_OUT, XNOR_1_3_NAND2_NUM396_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM396 (.ZN (XNOR_1_1_NAND2_NUM396_OUT), .A1 (N1252), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM396 (.ZN (XNOR_1_2_NAND2_NUM396_OUT), .A1 (GND), .A2 (N1253));
      NOR2_X1 XNOR_1_3_NAND2_NUM396 (.ZN (XNOR_1_3_NAND2_NUM396_OUT), .A1 (XNOR_1_1_NAND2_NUM396_OUT), .A2 (XNOR_1_2_NAND2_NUM396_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM396 (.ZN (N1304), .A1 (XNOR_1_3_NAND2_NUM396_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM397_OUT, XNOR_1_2_NAND2_NUM397_OUT, XNOR_1_3_NAND2_NUM397_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM397 (.ZN (XNOR_1_1_NAND2_NUM397_OUT), .A1 (N1254), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM397 (.ZN (XNOR_1_2_NAND2_NUM397_OUT), .A1 (GND), .A2 (N1255));
      NOR2_X1 XNOR_1_3_NAND2_NUM397 (.ZN (XNOR_1_3_NAND2_NUM397_OUT), .A1 (XNOR_1_1_NAND2_NUM397_OUT), .A2 (XNOR_1_2_NAND2_NUM397_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM397 (.ZN (N1305), .A1 (XNOR_1_3_NAND2_NUM397_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM398_OUT, XNOR_1_2_NAND2_NUM398_OUT, XNOR_1_3_NAND2_NUM398_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM398 (.ZN (XNOR_1_1_NAND2_NUM398_OUT), .A1 (N1256), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM398 (.ZN (XNOR_1_2_NAND2_NUM398_OUT), .A1 (GND), .A2 (N1257));
      NOR2_X1 XNOR_1_3_NAND2_NUM398 (.ZN (XNOR_1_3_NAND2_NUM398_OUT), .A1 (XNOR_1_1_NAND2_NUM398_OUT), .A2 (XNOR_1_2_NAND2_NUM398_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM398 (.ZN (N1306), .A1 (XNOR_1_3_NAND2_NUM398_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM399_OUT, XNOR_1_2_NAND2_NUM399_OUT, XNOR_1_3_NAND2_NUM399_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM399 (.ZN (XNOR_1_1_NAND2_NUM399_OUT), .A1 (N1258), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM399 (.ZN (XNOR_1_2_NAND2_NUM399_OUT), .A1 (GND), .A2 (N1259));
      NOR2_X1 XNOR_1_3_NAND2_NUM399 (.ZN (XNOR_1_3_NAND2_NUM399_OUT), .A1 (XNOR_1_1_NAND2_NUM399_OUT), .A2 (XNOR_1_2_NAND2_NUM399_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM399 (.ZN (N1307), .A1 (XNOR_1_3_NAND2_NUM399_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM400_OUT, XNOR_1_2_NAND2_NUM400_OUT, XNOR_1_3_NAND2_NUM400_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM400 (.ZN (XNOR_1_1_NAND2_NUM400_OUT), .A1 (N1260), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM400 (.ZN (XNOR_1_2_NAND2_NUM400_OUT), .A1 (GND), .A2 (N1261));
      NOR2_X1 XNOR_1_3_NAND2_NUM400 (.ZN (XNOR_1_3_NAND2_NUM400_OUT), .A1 (XNOR_1_1_NAND2_NUM400_OUT), .A2 (XNOR_1_2_NAND2_NUM400_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM400 (.ZN (N1308), .A1 (XNOR_1_3_NAND2_NUM400_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM401_OUT, XNOR_1_2_NAND2_NUM401_OUT, XNOR_1_3_NAND2_NUM401_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM401 (.ZN (XNOR_1_1_NAND2_NUM401_OUT), .A1 (N1262), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM401 (.ZN (XNOR_1_2_NAND2_NUM401_OUT), .A1 (GND), .A2 (N1263));
      NOR2_X1 XNOR_1_3_NAND2_NUM401 (.ZN (XNOR_1_3_NAND2_NUM401_OUT), .A1 (XNOR_1_1_NAND2_NUM401_OUT), .A2 (XNOR_1_2_NAND2_NUM401_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM401 (.ZN (N1309), .A1 (XNOR_1_3_NAND2_NUM401_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM402_OUT, XNOR_1_2_NAND2_NUM402_OUT, XNOR_1_3_NAND2_NUM402_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM402 (.ZN (XNOR_1_1_NAND2_NUM402_OUT), .A1 (N1264), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM402 (.ZN (XNOR_1_2_NAND2_NUM402_OUT), .A1 (GND), .A2 (N1265));
      NOR2_X1 XNOR_1_3_NAND2_NUM402 (.ZN (XNOR_1_3_NAND2_NUM402_OUT), .A1 (XNOR_1_1_NAND2_NUM402_OUT), .A2 (XNOR_1_2_NAND2_NUM402_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM402 (.ZN (N1310), .A1 (XNOR_1_3_NAND2_NUM402_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM403_OUT, XNOR_1_2_NAND2_NUM403_OUT, XNOR_1_3_NAND2_NUM403_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM403 (.ZN (XNOR_1_1_NAND2_NUM403_OUT), .A1 (N1266), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM403 (.ZN (XNOR_1_2_NAND2_NUM403_OUT), .A1 (GND), .A2 (N1267));
      NOR2_X1 XNOR_1_3_NAND2_NUM403 (.ZN (XNOR_1_3_NAND2_NUM403_OUT), .A1 (XNOR_1_1_NAND2_NUM403_OUT), .A2 (XNOR_1_2_NAND2_NUM403_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM403 (.ZN (N1311), .A1 (XNOR_1_3_NAND2_NUM403_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM404_OUT, XNOR_1_2_NAND2_NUM404_OUT, XNOR_1_3_NAND2_NUM404_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM404 (.ZN (XNOR_1_1_NAND2_NUM404_OUT), .A1 (N1268), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM404 (.ZN (XNOR_1_2_NAND2_NUM404_OUT), .A1 (GND), .A2 (N1269));
      NOR2_X1 XNOR_1_3_NAND2_NUM404 (.ZN (XNOR_1_3_NAND2_NUM404_OUT), .A1 (XNOR_1_1_NAND2_NUM404_OUT), .A2 (XNOR_1_2_NAND2_NUM404_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM404 (.ZN (N1312), .A1 (XNOR_1_3_NAND2_NUM404_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM405_OUT, XNOR_1_2_NAND2_NUM405_OUT, XNOR_1_3_NAND2_NUM405_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM405 (.ZN (XNOR_1_1_NAND2_NUM405_OUT), .A1 (N1270), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM405 (.ZN (XNOR_1_2_NAND2_NUM405_OUT), .A1 (GND), .A2 (N1271));
      NOR2_X1 XNOR_1_3_NAND2_NUM405 (.ZN (XNOR_1_3_NAND2_NUM405_OUT), .A1 (XNOR_1_1_NAND2_NUM405_OUT), .A2 (XNOR_1_2_NAND2_NUM405_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM405 (.ZN (N1313), .A1 (XNOR_1_3_NAND2_NUM405_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM406_OUT, XNOR_1_2_NAND2_NUM406_OUT, XNOR_1_3_NAND2_NUM406_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM406 (.ZN (XNOR_1_1_NAND2_NUM406_OUT), .A1 (N1272), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM406 (.ZN (XNOR_1_2_NAND2_NUM406_OUT), .A1 (GND), .A2 (N1273));
      NOR2_X1 XNOR_1_3_NAND2_NUM406 (.ZN (XNOR_1_3_NAND2_NUM406_OUT), .A1 (XNOR_1_1_NAND2_NUM406_OUT), .A2 (XNOR_1_2_NAND2_NUM406_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM406 (.ZN (N1314), .A1 (XNOR_1_3_NAND2_NUM406_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM407_OUT, XNOR_1_2_NAND2_NUM407_OUT, XNOR_1_3_NAND2_NUM407_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM407 (.ZN (XNOR_1_1_NAND2_NUM407_OUT), .A1 (N1274), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM407 (.ZN (XNOR_1_2_NAND2_NUM407_OUT), .A1 (GND), .A2 (N1275));
      NOR2_X1 XNOR_1_3_NAND2_NUM407 (.ZN (XNOR_1_3_NAND2_NUM407_OUT), .A1 (XNOR_1_1_NAND2_NUM407_OUT), .A2 (XNOR_1_2_NAND2_NUM407_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM407 (.ZN (N1315), .A1 (XNOR_1_3_NAND2_NUM407_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM408_OUT, XNOR_1_2_NAND2_NUM408_OUT, XNOR_1_3_NAND2_NUM408_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM408 (.ZN (XNOR_1_1_NAND2_NUM408_OUT), .A1 (N1276), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM408 (.ZN (XNOR_1_2_NAND2_NUM408_OUT), .A1 (GND), .A2 (N1277));
      NOR2_X1 XNOR_1_3_NAND2_NUM408 (.ZN (XNOR_1_3_NAND2_NUM408_OUT), .A1 (XNOR_1_1_NAND2_NUM408_OUT), .A2 (XNOR_1_2_NAND2_NUM408_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM408 (.ZN (N1316), .A1 (XNOR_1_3_NAND2_NUM408_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM409_OUT, XNOR_1_2_NAND2_NUM409_OUT, XNOR_1_3_NAND2_NUM409_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM409 (.ZN (XNOR_1_1_NAND2_NUM409_OUT), .A1 (N1278), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM409 (.ZN (XNOR_1_2_NAND2_NUM409_OUT), .A1 (GND), .A2 (N1279));
      NOR2_X1 XNOR_1_3_NAND2_NUM409 (.ZN (XNOR_1_3_NAND2_NUM409_OUT), .A1 (XNOR_1_1_NAND2_NUM409_OUT), .A2 (XNOR_1_2_NAND2_NUM409_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM409 (.ZN (N1317), .A1 (XNOR_1_3_NAND2_NUM409_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM410_OUT, XNOR_1_2_NAND2_NUM410_OUT, XNOR_1_3_NAND2_NUM410_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM410 (.ZN (XNOR_1_1_NAND2_NUM410_OUT), .A1 (N1280), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM410 (.ZN (XNOR_1_2_NAND2_NUM410_OUT), .A1 (GND), .A2 (N1281));
      NOR2_X1 XNOR_1_3_NAND2_NUM410 (.ZN (XNOR_1_3_NAND2_NUM410_OUT), .A1 (XNOR_1_1_NAND2_NUM410_OUT), .A2 (XNOR_1_2_NAND2_NUM410_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM410 (.ZN (N1318), .A1 (XNOR_1_3_NAND2_NUM410_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM411_OUT, XNOR_1_2_NAND2_NUM411_OUT, XNOR_1_3_NAND2_NUM411_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM411 (.ZN (XNOR_1_1_NAND2_NUM411_OUT), .A1 (N1282), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM411 (.ZN (XNOR_1_2_NAND2_NUM411_OUT), .A1 (GND), .A2 (N1283));
      NOR2_X1 XNOR_1_3_NAND2_NUM411 (.ZN (XNOR_1_3_NAND2_NUM411_OUT), .A1 (XNOR_1_1_NAND2_NUM411_OUT), .A2 (XNOR_1_2_NAND2_NUM411_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM411 (.ZN (N1319), .A1 (XNOR_1_3_NAND2_NUM411_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM412_OUT, XNOR_1_2_NAND2_NUM412_OUT, XNOR_1_3_NAND2_NUM412_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM412 (.ZN (XNOR_1_1_NAND2_NUM412_OUT), .A1 (N1284), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM412 (.ZN (XNOR_1_2_NAND2_NUM412_OUT), .A1 (GND), .A2 (N1285));
      NOR2_X1 XNOR_1_3_NAND2_NUM412 (.ZN (XNOR_1_3_NAND2_NUM412_OUT), .A1 (XNOR_1_1_NAND2_NUM412_OUT), .A2 (XNOR_1_2_NAND2_NUM412_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM412 (.ZN (N1320), .A1 (XNOR_1_3_NAND2_NUM412_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM413_OUT, XNOR_1_2_NAND2_NUM413_OUT, XNOR_1_3_NAND2_NUM413_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM413 (.ZN (XNOR_1_1_NAND2_NUM413_OUT), .A1 (N1286), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM413 (.ZN (XNOR_1_2_NAND2_NUM413_OUT), .A1 (GND), .A2 (N1287));
      NOR2_X1 XNOR_1_3_NAND2_NUM413 (.ZN (XNOR_1_3_NAND2_NUM413_OUT), .A1 (XNOR_1_1_NAND2_NUM413_OUT), .A2 (XNOR_1_2_NAND2_NUM413_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM413 (.ZN (N1321), .A1 (XNOR_1_3_NAND2_NUM413_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM414_OUT, XNOR_1_2_NAND2_NUM414_OUT, XNOR_1_3_NAND2_NUM414_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM414 (.ZN (XNOR_1_1_NAND2_NUM414_OUT), .A1 (N1288), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM414 (.ZN (XNOR_1_2_NAND2_NUM414_OUT), .A1 (GND), .A2 (N1289));
      NOR2_X1 XNOR_1_3_NAND2_NUM414 (.ZN (XNOR_1_3_NAND2_NUM414_OUT), .A1 (XNOR_1_1_NAND2_NUM414_OUT), .A2 (XNOR_1_2_NAND2_NUM414_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM414 (.ZN (N1322), .A1 (XNOR_1_3_NAND2_NUM414_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM415_OUT, XNOR_1_2_NAND2_NUM415_OUT, XNOR_1_3_NAND2_NUM415_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM415 (.ZN (XNOR_1_1_NAND2_NUM415_OUT), .A1 (N1290), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM415 (.ZN (XNOR_1_2_NAND2_NUM415_OUT), .A1 (GND), .A2 (N1291));
      NOR2_X1 XNOR_1_3_NAND2_NUM415 (.ZN (XNOR_1_3_NAND2_NUM415_OUT), .A1 (XNOR_1_1_NAND2_NUM415_OUT), .A2 (XNOR_1_2_NAND2_NUM415_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM415 (.ZN (N1323), .A1 (XNOR_1_3_NAND2_NUM415_OUT), .A2 (GND));
      wire XNOR_1_1_BUFF1_NUM0_OUT;
      NOR2_X1 XNOR_1_1_BUFF1_NUM0 (.ZN (XNOR_1_1_BUFF1_NUM0_OUT), .A1 (N1292), .A2 (GND));
      NOR2_X1 XNOR_1_2_BUFF1_NUM0 (.ZN (N1324), .A1 (XNOR_1_1_BUFF1_NUM0_OUT), .A2 (GND));
      wire XNOR_1_1_BUFF1_NUM1_OUT;
      NOR2_X1 XNOR_1_1_BUFF1_NUM1 (.ZN (XNOR_1_1_BUFF1_NUM1_OUT), .A1 (N1293), .A2 (GND));
      NOR2_X1 XNOR_1_2_BUFF1_NUM1 (.ZN (N1325), .A1 (XNOR_1_1_BUFF1_NUM1_OUT), .A2 (GND));
      wire XNOR_1_1_BUFF1_NUM2_OUT;
      NOR2_X1 XNOR_1_1_BUFF1_NUM2 (.ZN (XNOR_1_1_BUFF1_NUM2_OUT), .A1 (N1294), .A2 (GND));
      NOR2_X1 XNOR_1_2_BUFF1_NUM2 (.ZN (N1326), .A1 (XNOR_1_1_BUFF1_NUM2_OUT), .A2 (GND));
      wire XNOR_1_1_BUFF1_NUM3_OUT;
      NOR2_X1 XNOR_1_1_BUFF1_NUM3 (.ZN (XNOR_1_1_BUFF1_NUM3_OUT), .A1 (N1295), .A2 (GND));
      NOR2_X1 XNOR_1_2_BUFF1_NUM3 (.ZN (N1327), .A1 (XNOR_1_1_BUFF1_NUM3_OUT), .A2 (GND));
      wire XNOR_1_1_BUFF1_NUM4_OUT;
      NOR2_X1 XNOR_1_1_BUFF1_NUM4 (.ZN (XNOR_1_1_BUFF1_NUM4_OUT), .A1 (N1296), .A2 (GND));
      NOR2_X1 XNOR_1_2_BUFF1_NUM4 (.ZN (N1328), .A1 (XNOR_1_1_BUFF1_NUM4_OUT), .A2 (GND));
      wire XNOR_1_1_BUFF1_NUM5_OUT;
      NOR2_X1 XNOR_1_1_BUFF1_NUM5 (.ZN (XNOR_1_1_BUFF1_NUM5_OUT), .A1 (N1297), .A2 (GND));
      NOR2_X1 XNOR_1_2_BUFF1_NUM5 (.ZN (N1329), .A1 (XNOR_1_1_BUFF1_NUM5_OUT), .A2 (GND));
      wire XNOR_1_1_BUFF1_NUM6_OUT;
      NOR2_X1 XNOR_1_1_BUFF1_NUM6 (.ZN (XNOR_1_1_BUFF1_NUM6_OUT), .A1 (N1298), .A2 (GND));
      NOR2_X1 XNOR_1_2_BUFF1_NUM6 (.ZN (N1330), .A1 (XNOR_1_1_BUFF1_NUM6_OUT), .A2 (GND));
      wire XNOR_1_1_BUFF1_NUM7_OUT;
      NOR2_X1 XNOR_1_1_BUFF1_NUM7 (.ZN (XNOR_1_1_BUFF1_NUM7_OUT), .A1 (N1299), .A2 (GND));
      NOR2_X1 XNOR_1_2_BUFF1_NUM7 (.ZN (N1331), .A1 (XNOR_1_1_BUFF1_NUM7_OUT), .A2 (GND));
      wire XNOR_1_1_BUFF1_NUM8_OUT;
      NOR2_X1 XNOR_1_1_BUFF1_NUM8 (.ZN (XNOR_1_1_BUFF1_NUM8_OUT), .A1 (N1300), .A2 (GND));
      NOR2_X1 XNOR_1_2_BUFF1_NUM8 (.ZN (N1332), .A1 (XNOR_1_1_BUFF1_NUM8_OUT), .A2 (GND));
      wire XNOR_1_1_BUFF1_NUM9_OUT;
      NOR2_X1 XNOR_1_1_BUFF1_NUM9 (.ZN (XNOR_1_1_BUFF1_NUM9_OUT), .A1 (N1301), .A2 (GND));
      NOR2_X1 XNOR_1_2_BUFF1_NUM9 (.ZN (N1333), .A1 (XNOR_1_1_BUFF1_NUM9_OUT), .A2 (GND));
      wire XNOR_1_1_BUFF1_NUM10_OUT;
      NOR2_X1 XNOR_1_1_BUFF1_NUM10 (.ZN (XNOR_1_1_BUFF1_NUM10_OUT), .A1 (N1302), .A2 (GND));
      NOR2_X1 XNOR_1_2_BUFF1_NUM10 (.ZN (N1334), .A1 (XNOR_1_1_BUFF1_NUM10_OUT), .A2 (GND));
      wire XNOR_1_1_BUFF1_NUM11_OUT;
      NOR2_X1 XNOR_1_1_BUFF1_NUM11 (.ZN (XNOR_1_1_BUFF1_NUM11_OUT), .A1 (N1303), .A2 (GND));
      NOR2_X1 XNOR_1_2_BUFF1_NUM11 (.ZN (N1335), .A1 (XNOR_1_1_BUFF1_NUM11_OUT), .A2 (GND));
      wire XNOR_1_1_BUFF1_NUM12_OUT;
      NOR2_X1 XNOR_1_1_BUFF1_NUM12 (.ZN (XNOR_1_1_BUFF1_NUM12_OUT), .A1 (N1304), .A2 (GND));
      NOR2_X1 XNOR_1_2_BUFF1_NUM12 (.ZN (N1336), .A1 (XNOR_1_1_BUFF1_NUM12_OUT), .A2 (GND));
      wire XNOR_1_1_BUFF1_NUM13_OUT;
      NOR2_X1 XNOR_1_1_BUFF1_NUM13 (.ZN (XNOR_1_1_BUFF1_NUM13_OUT), .A1 (N1305), .A2 (GND));
      NOR2_X1 XNOR_1_2_BUFF1_NUM13 (.ZN (N1337), .A1 (XNOR_1_1_BUFF1_NUM13_OUT), .A2 (GND));
      wire XNOR_1_1_BUFF1_NUM14_OUT;
      NOR2_X1 XNOR_1_1_BUFF1_NUM14 (.ZN (XNOR_1_1_BUFF1_NUM14_OUT), .A1 (N1306), .A2 (GND));
      NOR2_X1 XNOR_1_2_BUFF1_NUM14 (.ZN (N1338), .A1 (XNOR_1_1_BUFF1_NUM14_OUT), .A2 (GND));
      wire XNOR_1_1_BUFF1_NUM15_OUT;
      NOR2_X1 XNOR_1_1_BUFF1_NUM15 (.ZN (XNOR_1_1_BUFF1_NUM15_OUT), .A1 (N1307), .A2 (GND));
      NOR2_X1 XNOR_1_2_BUFF1_NUM15 (.ZN (N1339), .A1 (XNOR_1_1_BUFF1_NUM15_OUT), .A2 (GND));
      wire XNOR_1_1_BUFF1_NUM16_OUT;
      NOR2_X1 XNOR_1_1_BUFF1_NUM16 (.ZN (XNOR_1_1_BUFF1_NUM16_OUT), .A1 (N1308), .A2 (GND));
      NOR2_X1 XNOR_1_2_BUFF1_NUM16 (.ZN (N1340), .A1 (XNOR_1_1_BUFF1_NUM16_OUT), .A2 (GND));
      wire XNOR_1_1_BUFF1_NUM17_OUT;
      NOR2_X1 XNOR_1_1_BUFF1_NUM17 (.ZN (XNOR_1_1_BUFF1_NUM17_OUT), .A1 (N1309), .A2 (GND));
      NOR2_X1 XNOR_1_2_BUFF1_NUM17 (.ZN (N1341), .A1 (XNOR_1_1_BUFF1_NUM17_OUT), .A2 (GND));
      wire XNOR_1_1_BUFF1_NUM18_OUT;
      NOR2_X1 XNOR_1_1_BUFF1_NUM18 (.ZN (XNOR_1_1_BUFF1_NUM18_OUT), .A1 (N1310), .A2 (GND));
      NOR2_X1 XNOR_1_2_BUFF1_NUM18 (.ZN (N1342), .A1 (XNOR_1_1_BUFF1_NUM18_OUT), .A2 (GND));
      wire XNOR_1_1_BUFF1_NUM19_OUT;
      NOR2_X1 XNOR_1_1_BUFF1_NUM19 (.ZN (XNOR_1_1_BUFF1_NUM19_OUT), .A1 (N1311), .A2 (GND));
      NOR2_X1 XNOR_1_2_BUFF1_NUM19 (.ZN (N1343), .A1 (XNOR_1_1_BUFF1_NUM19_OUT), .A2 (GND));
      wire XNOR_1_1_BUFF1_NUM20_OUT;
      NOR2_X1 XNOR_1_1_BUFF1_NUM20 (.ZN (XNOR_1_1_BUFF1_NUM20_OUT), .A1 (N1312), .A2 (GND));
      NOR2_X1 XNOR_1_2_BUFF1_NUM20 (.ZN (N1344), .A1 (XNOR_1_1_BUFF1_NUM20_OUT), .A2 (GND));
      wire XNOR_1_1_BUFF1_NUM21_OUT;
      NOR2_X1 XNOR_1_1_BUFF1_NUM21 (.ZN (XNOR_1_1_BUFF1_NUM21_OUT), .A1 (N1313), .A2 (GND));
      NOR2_X1 XNOR_1_2_BUFF1_NUM21 (.ZN (N1345), .A1 (XNOR_1_1_BUFF1_NUM21_OUT), .A2 (GND));
      wire XNOR_1_1_BUFF1_NUM22_OUT;
      NOR2_X1 XNOR_1_1_BUFF1_NUM22 (.ZN (XNOR_1_1_BUFF1_NUM22_OUT), .A1 (N1314), .A2 (GND));
      NOR2_X1 XNOR_1_2_BUFF1_NUM22 (.ZN (N1346), .A1 (XNOR_1_1_BUFF1_NUM22_OUT), .A2 (GND));
      wire XNOR_1_1_BUFF1_NUM23_OUT;
      NOR2_X1 XNOR_1_1_BUFF1_NUM23 (.ZN (XNOR_1_1_BUFF1_NUM23_OUT), .A1 (N1315), .A2 (GND));
      NOR2_X1 XNOR_1_2_BUFF1_NUM23 (.ZN (N1347), .A1 (XNOR_1_1_BUFF1_NUM23_OUT), .A2 (GND));
      wire XNOR_1_1_BUFF1_NUM24_OUT;
      NOR2_X1 XNOR_1_1_BUFF1_NUM24 (.ZN (XNOR_1_1_BUFF1_NUM24_OUT), .A1 (N1316), .A2 (GND));
      NOR2_X1 XNOR_1_2_BUFF1_NUM24 (.ZN (N1348), .A1 (XNOR_1_1_BUFF1_NUM24_OUT), .A2 (GND));
      wire XNOR_1_1_BUFF1_NUM25_OUT;
      NOR2_X1 XNOR_1_1_BUFF1_NUM25 (.ZN (XNOR_1_1_BUFF1_NUM25_OUT), .A1 (N1317), .A2 (GND));
      NOR2_X1 XNOR_1_2_BUFF1_NUM25 (.ZN (N1349), .A1 (XNOR_1_1_BUFF1_NUM25_OUT), .A2 (GND));
      wire XNOR_1_1_BUFF1_NUM26_OUT;
      NOR2_X1 XNOR_1_1_BUFF1_NUM26 (.ZN (XNOR_1_1_BUFF1_NUM26_OUT), .A1 (N1318), .A2 (GND));
      NOR2_X1 XNOR_1_2_BUFF1_NUM26 (.ZN (N1350), .A1 (XNOR_1_1_BUFF1_NUM26_OUT), .A2 (GND));
      wire XNOR_1_1_BUFF1_NUM27_OUT;
      NOR2_X1 XNOR_1_1_BUFF1_NUM27 (.ZN (XNOR_1_1_BUFF1_NUM27_OUT), .A1 (N1319), .A2 (GND));
      NOR2_X1 XNOR_1_2_BUFF1_NUM27 (.ZN (N1351), .A1 (XNOR_1_1_BUFF1_NUM27_OUT), .A2 (GND));
      wire XNOR_1_1_BUFF1_NUM28_OUT;
      NOR2_X1 XNOR_1_1_BUFF1_NUM28 (.ZN (XNOR_1_1_BUFF1_NUM28_OUT), .A1 (N1320), .A2 (GND));
      NOR2_X1 XNOR_1_2_BUFF1_NUM28 (.ZN (N1352), .A1 (XNOR_1_1_BUFF1_NUM28_OUT), .A2 (GND));
      wire XNOR_1_1_BUFF1_NUM29_OUT;
      NOR2_X1 XNOR_1_1_BUFF1_NUM29 (.ZN (XNOR_1_1_BUFF1_NUM29_OUT), .A1 (N1321), .A2 (GND));
      NOR2_X1 XNOR_1_2_BUFF1_NUM29 (.ZN (N1353), .A1 (XNOR_1_1_BUFF1_NUM29_OUT), .A2 (GND));
      wire XNOR_1_1_BUFF1_NUM30_OUT;
      NOR2_X1 XNOR_1_1_BUFF1_NUM30 (.ZN (XNOR_1_1_BUFF1_NUM30_OUT), .A1 (N1322), .A2 (GND));
      NOR2_X1 XNOR_1_2_BUFF1_NUM30 (.ZN (N1354), .A1 (XNOR_1_1_BUFF1_NUM30_OUT), .A2 (GND));
      wire XNOR_1_1_BUFF1_NUM31_OUT;
      NOR2_X1 XNOR_1_1_BUFF1_NUM31 (.ZN (XNOR_1_1_BUFF1_NUM31_OUT), .A1 (N1323), .A2 (GND));
      NOR2_X1 XNOR_1_2_BUFF1_NUM31 (.ZN (N1355), .A1 (XNOR_1_1_BUFF1_NUM31_OUT), .A2 (GND));


      wire XNOR_1_1_N1324_TERMINATION_OUT, XNOR_1_2_N1324_TERMINATION_OUT;
      NOR2_X1 XNOR_1_1_N1324_TERMINATION (.ZN (XNOR_1_1_N1324_TERMINATION_OUT), .A1 (N1324), .A2 (GND));
      NOR2_X1 XNOR_1_2_N1324_TERMINATION (.ZN (N1324_TERMINATION), .A1 (XNOR_1_1_N1324_TERMINATION_OUT), .A2 (XNOR_1_2_N1324_TERMINATION_OUT));

      wire XNOR_1_1_N1325_TERMINATION_OUT, XNOR_1_2_N1325_TERMINATION_OUT;
      NOR2_X1 XNOR_1_1_N1325_TERMINATION (.ZN (XNOR_1_1_N1325_TERMINATION_OUT), .A1 (N1325), .A2 (GND));
      NOR2_X1 XNOR_1_2_N1325_TERMINATION (.ZN (N1325_TERMINATION), .A1 (XNOR_1_1_N1325_TERMINATION_OUT), .A2 (XNOR_1_2_N1325_TERMINATION_OUT));

      wire XNOR_1_1_N1326_TERMINATION_OUT, XNOR_1_2_N1326_TERMINATION_OUT;
      NOR2_X1 XNOR_1_1_N1326_TERMINATION (.ZN (XNOR_1_1_N1326_TERMINATION_OUT), .A1 (N1326), .A2 (GND));
      NOR2_X1 XNOR_1_2_N1326_TERMINATION (.ZN (N1326_TERMINATION), .A1 (XNOR_1_1_N1326_TERMINATION_OUT), .A2 (XNOR_1_2_N1326_TERMINATION_OUT));

      wire XNOR_1_1_N1327_TERMINATION_OUT, XNOR_1_2_N1327_TERMINATION_OUT;
      NOR2_X1 XNOR_1_1_N1327_TERMINATION (.ZN (XNOR_1_1_N1327_TERMINATION_OUT), .A1 (N1327), .A2 (GND));
      NOR2_X1 XNOR_1_2_N1327_TERMINATION (.ZN (N1327_TERMINATION), .A1 (XNOR_1_1_N1327_TERMINATION_OUT), .A2 (XNOR_1_2_N1327_TERMINATION_OUT));

      wire XNOR_1_1_N1328_TERMINATION_OUT, XNOR_1_2_N1328_TERMINATION_OUT;
      NOR2_X1 XNOR_1_1_N1328_TERMINATION (.ZN (XNOR_1_1_N1328_TERMINATION_OUT), .A1 (N1328), .A2 (GND));
      NOR2_X1 XNOR_1_2_N1328_TERMINATION (.ZN (N1328_TERMINATION), .A1 (XNOR_1_1_N1328_TERMINATION_OUT), .A2 (XNOR_1_2_N1328_TERMINATION_OUT));

      wire XNOR_1_1_N1329_TERMINATION_OUT, XNOR_1_2_N1329_TERMINATION_OUT;
      NOR2_X1 XNOR_1_1_N1329_TERMINATION (.ZN (XNOR_1_1_N1329_TERMINATION_OUT), .A1 (N1329), .A2 (GND));
      NOR2_X1 XNOR_1_2_N1329_TERMINATION (.ZN (N1329_TERMINATION), .A1 (XNOR_1_1_N1329_TERMINATION_OUT), .A2 (XNOR_1_2_N1329_TERMINATION_OUT));

      wire XNOR_1_1_N1330_TERMINATION_OUT, XNOR_1_2_N1330_TERMINATION_OUT;
      NOR2_X1 XNOR_1_1_N1330_TERMINATION (.ZN (XNOR_1_1_N1330_TERMINATION_OUT), .A1 (N1330), .A2 (GND));
      NOR2_X1 XNOR_1_2_N1330_TERMINATION (.ZN (N1330_TERMINATION), .A1 (XNOR_1_1_N1330_TERMINATION_OUT), .A2 (XNOR_1_2_N1330_TERMINATION_OUT));

      wire XNOR_1_1_N1331_TERMINATION_OUT, XNOR_1_2_N1331_TERMINATION_OUT;
      NOR2_X1 XNOR_1_1_N1331_TERMINATION (.ZN (XNOR_1_1_N1331_TERMINATION_OUT), .A1 (N1331), .A2 (GND));
      NOR2_X1 XNOR_1_2_N1331_TERMINATION (.ZN (N1331_TERMINATION), .A1 (XNOR_1_1_N1331_TERMINATION_OUT), .A2 (XNOR_1_2_N1331_TERMINATION_OUT));

      wire XNOR_1_1_N1332_TERMINATION_OUT, XNOR_1_2_N1332_TERMINATION_OUT;
      NOR2_X1 XNOR_1_1_N1332_TERMINATION (.ZN (XNOR_1_1_N1332_TERMINATION_OUT), .A1 (N1332), .A2 (GND));
      NOR2_X1 XNOR_1_2_N1332_TERMINATION (.ZN (N1332_TERMINATION), .A1 (XNOR_1_1_N1332_TERMINATION_OUT), .A2 (XNOR_1_2_N1332_TERMINATION_OUT));

      wire XNOR_1_1_N1333_TERMINATION_OUT, XNOR_1_2_N1333_TERMINATION_OUT;
      NOR2_X1 XNOR_1_1_N1333_TERMINATION (.ZN (XNOR_1_1_N1333_TERMINATION_OUT), .A1 (N1333), .A2 (GND));
      NOR2_X1 XNOR_1_2_N1333_TERMINATION (.ZN (N1333_TERMINATION), .A1 (XNOR_1_1_N1333_TERMINATION_OUT), .A2 (XNOR_1_2_N1333_TERMINATION_OUT));

      wire XNOR_1_1_N1334_TERMINATION_OUT, XNOR_1_2_N1334_TERMINATION_OUT;
      NOR2_X1 XNOR_1_1_N1334_TERMINATION (.ZN (XNOR_1_1_N1334_TERMINATION_OUT), .A1 (N1334), .A2 (GND));
      NOR2_X1 XNOR_1_2_N1334_TERMINATION (.ZN (N1334_TERMINATION), .A1 (XNOR_1_1_N1334_TERMINATION_OUT), .A2 (XNOR_1_2_N1334_TERMINATION_OUT));

      wire XNOR_1_1_N1335_TERMINATION_OUT, XNOR_1_2_N1335_TERMINATION_OUT;
      NOR2_X1 XNOR_1_1_N1335_TERMINATION (.ZN (XNOR_1_1_N1335_TERMINATION_OUT), .A1 (N1335), .A2 (GND));
      NOR2_X1 XNOR_1_2_N1335_TERMINATION (.ZN (N1335_TERMINATION), .A1 (XNOR_1_1_N1335_TERMINATION_OUT), .A2 (XNOR_1_2_N1335_TERMINATION_OUT));

      wire XNOR_1_1_N1336_TERMINATION_OUT, XNOR_1_2_N1336_TERMINATION_OUT;
      NOR2_X1 XNOR_1_1_N1336_TERMINATION (.ZN (XNOR_1_1_N1336_TERMINATION_OUT), .A1 (N1336), .A2 (GND));
      NOR2_X1 XNOR_1_2_N1336_TERMINATION (.ZN (N1336_TERMINATION), .A1 (XNOR_1_1_N1336_TERMINATION_OUT), .A2 (XNOR_1_2_N1336_TERMINATION_OUT));

      wire XNOR_1_1_N1337_TERMINATION_OUT, XNOR_1_2_N1337_TERMINATION_OUT;
      NOR2_X1 XNOR_1_1_N1337_TERMINATION (.ZN (XNOR_1_1_N1337_TERMINATION_OUT), .A1 (N1337), .A2 (GND));
      NOR2_X1 XNOR_1_2_N1337_TERMINATION (.ZN (N1337_TERMINATION), .A1 (XNOR_1_1_N1337_TERMINATION_OUT), .A2 (XNOR_1_2_N1337_TERMINATION_OUT));

      wire XNOR_1_1_N1338_TERMINATION_OUT, XNOR_1_2_N1338_TERMINATION_OUT;
      NOR2_X1 XNOR_1_1_N1338_TERMINATION (.ZN (XNOR_1_1_N1338_TERMINATION_OUT), .A1 (N1338), .A2 (GND));
      NOR2_X1 XNOR_1_2_N1338_TERMINATION (.ZN (N1338_TERMINATION), .A1 (XNOR_1_1_N1338_TERMINATION_OUT), .A2 (XNOR_1_2_N1338_TERMINATION_OUT));

      wire XNOR_1_1_N1339_TERMINATION_OUT, XNOR_1_2_N1339_TERMINATION_OUT;
      NOR2_X1 XNOR_1_1_N1339_TERMINATION (.ZN (XNOR_1_1_N1339_TERMINATION_OUT), .A1 (N1339), .A2 (GND));
      NOR2_X1 XNOR_1_2_N1339_TERMINATION (.ZN (N1339_TERMINATION), .A1 (XNOR_1_1_N1339_TERMINATION_OUT), .A2 (XNOR_1_2_N1339_TERMINATION_OUT));

      wire XNOR_1_1_N1340_TERMINATION_OUT, XNOR_1_2_N1340_TERMINATION_OUT;
      NOR2_X1 XNOR_1_1_N1340_TERMINATION (.ZN (XNOR_1_1_N1340_TERMINATION_OUT), .A1 (N1340), .A2 (GND));
      NOR2_X1 XNOR_1_2_N1340_TERMINATION (.ZN (N1340_TERMINATION), .A1 (XNOR_1_1_N1340_TERMINATION_OUT), .A2 (XNOR_1_2_N1340_TERMINATION_OUT));

      wire XNOR_1_1_N1341_TERMINATION_OUT, XNOR_1_2_N1341_TERMINATION_OUT;
      NOR2_X1 XNOR_1_1_N1341_TERMINATION (.ZN (XNOR_1_1_N1341_TERMINATION_OUT), .A1 (N1341), .A2 (GND));
      NOR2_X1 XNOR_1_2_N1341_TERMINATION (.ZN (N1341_TERMINATION), .A1 (XNOR_1_1_N1341_TERMINATION_OUT), .A2 (XNOR_1_2_N1341_TERMINATION_OUT));

      wire XNOR_1_1_N1342_TERMINATION_OUT, XNOR_1_2_N1342_TERMINATION_OUT;
      NOR2_X1 XNOR_1_1_N1342_TERMINATION (.ZN (XNOR_1_1_N1342_TERMINATION_OUT), .A1 (N1342), .A2 (GND));
      NOR2_X1 XNOR_1_2_N1342_TERMINATION (.ZN (N1342_TERMINATION), .A1 (XNOR_1_1_N1342_TERMINATION_OUT), .A2 (XNOR_1_2_N1342_TERMINATION_OUT));

      wire XNOR_1_1_N1343_TERMINATION_OUT, XNOR_1_2_N1343_TERMINATION_OUT;
      NOR2_X1 XNOR_1_1_N1343_TERMINATION (.ZN (XNOR_1_1_N1343_TERMINATION_OUT), .A1 (N1343), .A2 (GND));
      NOR2_X1 XNOR_1_2_N1343_TERMINATION (.ZN (N1343_TERMINATION), .A1 (XNOR_1_1_N1343_TERMINATION_OUT), .A2 (XNOR_1_2_N1343_TERMINATION_OUT));

      wire XNOR_1_1_N1344_TERMINATION_OUT, XNOR_1_2_N1344_TERMINATION_OUT;
      NOR2_X1 XNOR_1_1_N1344_TERMINATION (.ZN (XNOR_1_1_N1344_TERMINATION_OUT), .A1 (N1344), .A2 (GND));
      NOR2_X1 XNOR_1_2_N1344_TERMINATION (.ZN (N1344_TERMINATION), .A1 (XNOR_1_1_N1344_TERMINATION_OUT), .A2 (XNOR_1_2_N1344_TERMINATION_OUT));

      wire XNOR_1_1_N1345_TERMINATION_OUT, XNOR_1_2_N1345_TERMINATION_OUT;
      NOR2_X1 XNOR_1_1_N1345_TERMINATION (.ZN (XNOR_1_1_N1345_TERMINATION_OUT), .A1 (N1345), .A2 (GND));
      NOR2_X1 XNOR_1_2_N1345_TERMINATION (.ZN (N1345_TERMINATION), .A1 (XNOR_1_1_N1345_TERMINATION_OUT), .A2 (XNOR_1_2_N1345_TERMINATION_OUT));

      wire XNOR_1_1_N1346_TERMINATION_OUT, XNOR_1_2_N1346_TERMINATION_OUT;
      NOR2_X1 XNOR_1_1_N1346_TERMINATION (.ZN (XNOR_1_1_N1346_TERMINATION_OUT), .A1 (N1346), .A2 (GND));
      NOR2_X1 XNOR_1_2_N1346_TERMINATION (.ZN (N1346_TERMINATION), .A1 (XNOR_1_1_N1346_TERMINATION_OUT), .A2 (XNOR_1_2_N1346_TERMINATION_OUT));

      wire XNOR_1_1_N1347_TERMINATION_OUT, XNOR_1_2_N1347_TERMINATION_OUT;
      NOR2_X1 XNOR_1_1_N1347_TERMINATION (.ZN (XNOR_1_1_N1347_TERMINATION_OUT), .A1 (N1347), .A2 (GND));
      NOR2_X1 XNOR_1_2_N1347_TERMINATION (.ZN (N1347_TERMINATION), .A1 (XNOR_1_1_N1347_TERMINATION_OUT), .A2 (XNOR_1_2_N1347_TERMINATION_OUT));

      wire XNOR_1_1_N1348_TERMINATION_OUT, XNOR_1_2_N1348_TERMINATION_OUT;
      NOR2_X1 XNOR_1_1_N1348_TERMINATION (.ZN (XNOR_1_1_N1348_TERMINATION_OUT), .A1 (N1348), .A2 (GND));
      NOR2_X1 XNOR_1_2_N1348_TERMINATION (.ZN (N1348_TERMINATION), .A1 (XNOR_1_1_N1348_TERMINATION_OUT), .A2 (XNOR_1_2_N1348_TERMINATION_OUT));

      wire XNOR_1_1_N1349_TERMINATION_OUT, XNOR_1_2_N1349_TERMINATION_OUT;
      NOR2_X1 XNOR_1_1_N1349_TERMINATION (.ZN (XNOR_1_1_N1349_TERMINATION_OUT), .A1 (N1349), .A2 (GND));
      NOR2_X1 XNOR_1_2_N1349_TERMINATION (.ZN (N1349_TERMINATION), .A1 (XNOR_1_1_N1349_TERMINATION_OUT), .A2 (XNOR_1_2_N1349_TERMINATION_OUT));

      wire XNOR_1_1_N1350_TERMINATION_OUT, XNOR_1_2_N1350_TERMINATION_OUT;
      NOR2_X1 XNOR_1_1_N1350_TERMINATION (.ZN (XNOR_1_1_N1350_TERMINATION_OUT), .A1 (N1350), .A2 (GND));
      NOR2_X1 XNOR_1_2_N1350_TERMINATION (.ZN (N1350_TERMINATION), .A1 (XNOR_1_1_N1350_TERMINATION_OUT), .A2 (XNOR_1_2_N1350_TERMINATION_OUT));

      wire XNOR_1_1_N1351_TERMINATION_OUT, XNOR_1_2_N1351_TERMINATION_OUT;
      NOR2_X1 XNOR_1_1_N1351_TERMINATION (.ZN (XNOR_1_1_N1351_TERMINATION_OUT), .A1 (N1351), .A2 (GND));
      NOR2_X1 XNOR_1_2_N1351_TERMINATION (.ZN (N1351_TERMINATION), .A1 (XNOR_1_1_N1351_TERMINATION_OUT), .A2 (XNOR_1_2_N1351_TERMINATION_OUT));

      wire XNOR_1_1_N1352_TERMINATION_OUT, XNOR_1_2_N1352_TERMINATION_OUT;
      NOR2_X1 XNOR_1_1_N1352_TERMINATION (.ZN (XNOR_1_1_N1352_TERMINATION_OUT), .A1 (N1352), .A2 (GND));
      NOR2_X1 XNOR_1_2_N1352_TERMINATION (.ZN (N1352_TERMINATION), .A1 (XNOR_1_1_N1352_TERMINATION_OUT), .A2 (XNOR_1_2_N1352_TERMINATION_OUT));

      wire XNOR_1_1_N1353_TERMINATION_OUT, XNOR_1_2_N1353_TERMINATION_OUT;
      NOR2_X1 XNOR_1_1_N1353_TERMINATION (.ZN (XNOR_1_1_N1353_TERMINATION_OUT), .A1 (N1353), .A2 (GND));
      NOR2_X1 XNOR_1_2_N1353_TERMINATION (.ZN (N1353_TERMINATION), .A1 (XNOR_1_1_N1353_TERMINATION_OUT), .A2 (XNOR_1_2_N1353_TERMINATION_OUT));

      wire XNOR_1_1_N1354_TERMINATION_OUT, XNOR_1_2_N1354_TERMINATION_OUT;
      NOR2_X1 XNOR_1_1_N1354_TERMINATION (.ZN (XNOR_1_1_N1354_TERMINATION_OUT), .A1 (N1354), .A2 (GND));
      NOR2_X1 XNOR_1_2_N1354_TERMINATION (.ZN (N1354_TERMINATION), .A1 (XNOR_1_1_N1354_TERMINATION_OUT), .A2 (XNOR_1_2_N1354_TERMINATION_OUT));

      wire XNOR_1_1_N1355_TERMINATION_OUT, XNOR_1_2_N1355_TERMINATION_OUT;
      NOR2_X1 XNOR_1_1_N1355_TERMINATION (.ZN (XNOR_1_1_N1355_TERMINATION_OUT), .A1 (N1355), .A2 (GND));
      NOR2_X1 XNOR_1_2_N1355_TERMINATION (.ZN (N1355_TERMINATION), .A1 (XNOR_1_1_N1355_TERMINATION_OUT), .A2 (XNOR_1_2_N1355_TERMINATION_OUT));





endmodule
* circuit: nor_funnel
simulator lang=spice

*.PARAM pw=<sed>pw<sed>as
.PARAM supp=0.8V slope=0.1fs
.PARAM t_init0=0.1ns t_init1=0.174ns
.PARAM baseVal=0V peakVal=0.8V tend=1.0ns


.LIB /home/s11777724/involution_tool_library_files/backend/spice/fet.inc CMG

* main circuit
.INCLUDE /home/s11777724/involution_tool_library_files/backend/spice/cell/NOR2_X1.sp
.INCLUDE /home/s11777724/involution_tool_library_files/backend/spice/cell/INV_X1.sp

**** SPECTRE Back Annotation
.option spef='/home/s11777724/JS/idm_evaluation/nor_funnel/place_and_route/nor_funnel_generic_parasitics.spef'
****

.TEMP 25
.OPTION
+ INGOLD=2
+ PARHIER=LOCAL
*+ POST=CSDF
+ PROBE
+ BRIEF
+ ACCURATE
+ ABSVAR=0.0001
+ DVDT=2
+ RELTOL=1e-11
*+ DELMAX=100fs
+ dc_pivot_check=yes

* vdd
VDD VDD GND 0.8v

* circuit under test

XINV_STAGE_0 STAGE_1_OUT STAGE_0_INTERNAL VDD VDD GND GND INV_X1
XNOR_STAGE_0 STAGE_29_OUT STAGE_0_INTERNAL STAGE_0_OUT VDD VDD GND GND NOR2_X1

XINV_STAGE_1 STAGE_2_OUT STAGE_1_INTERNAL VDD VDD GND GND INV_X1
XNOR_STAGE_1 STAGE_0_OUT STAGE_1_INTERNAL STAGE_1_OUT VDD VDD GND GND NOR2_X1

XINV_STAGE_2 STAGE_3_OUT STAGE_2_INTERNAL VDD VDD GND GND INV_X1
XNOR_STAGE_2 STAGE_1_OUT STAGE_2_INTERNAL STAGE_2_OUT VDD VDD GND GND NOR2_X1

XINV_STAGE_3 STAGE_4_OUT STAGE_3_INTERNAL VDD VDD GND GND INV_X1
XNOR_STAGE_3 STAGE_2_OUT STAGE_3_INTERNAL STAGE_3_OUT VDD VDD GND GND NOR2_X1

XINV_STAGE_4 STAGE_5_OUT STAGE_4_INTERNAL VDD VDD GND GND INV_X1
XNOR_STAGE_4 STAGE_3_OUT STAGE_4_INTERNAL STAGE_4_OUT VDD VDD GND GND NOR2_X1

XINV_STAGE_5 STAGE_6_OUT STAGE_5_INTERNAL VDD VDD GND GND INV_X1
XNOR_STAGE_5 STAGE_4_OUT STAGE_5_INTERNAL STAGE_5_OUT VDD VDD GND GND NOR2_X1

XINV_STAGE_6 STAGE_7_OUT STAGE_6_INTERNAL VDD VDD GND GND INV_X1
XNOR_STAGE_6 STAGE_5_OUT STAGE_6_INTERNAL STAGE_6_OUT VDD VDD GND GND NOR2_X1

XINV_STAGE_7 STAGE_8_OUT STAGE_7_INTERNAL VDD VDD GND GND INV_X1
XNOR_STAGE_7 STAGE_6_OUT STAGE_7_INTERNAL STAGE_7_OUT VDD VDD GND GND NOR2_X1

XINV_STAGE_8 STAGE_9_OUT STAGE_8_INTERNAL VDD VDD GND GND INV_X1
XNOR_STAGE_8 STAGE_7_OUT STAGE_8_INTERNAL STAGE_8_OUT VDD VDD GND GND NOR2_X1

XINV_STAGE_9 STAGE_10_OUT STAGE_9_INTERNAL VDD VDD GND GND INV_X1
XNOR_STAGE_9 STAGE_8_OUT STAGE_9_INTERNAL STAGE_9_OUT VDD VDD GND GND NOR2_X1

XINV_STAGE_10 STAGE_11_OUT STAGE_10_INTERNAL VDD VDD GND GND INV_X1
XNOR_STAGE_10 STAGE_9_OUT STAGE_10_INTERNAL STAGE_10_OUT VDD VDD GND GND NOR2_X1

XINV_STAGE_11 STAGE_12_OUT STAGE_11_INTERNAL VDD VDD GND GND INV_X1
XNOR_STAGE_11 STAGE_10_OUT STAGE_11_INTERNAL STAGE_11_OUT VDD VDD GND GND NOR2_X1

XINV_STAGE_12 STAGE_13_OUT STAGE_12_INTERNAL VDD VDD GND GND INV_X1
XNOR_STAGE_12 STAGE_11_OUT STAGE_12_INTERNAL STAGE_12_OUT VDD VDD GND GND NOR2_X1

XINV_STAGE_13 STAGE_14_OUT STAGE_13_INTERNAL VDD VDD GND GND INV_X1
XNOR_STAGE_13 STAGE_12_OUT STAGE_13_INTERNAL STAGE_13_OUT VDD VDD GND GND NOR2_X1

XINV_STAGE_14 STAGE_15_OUT STAGE_14_INTERNAL VDD VDD GND GND INV_X1
XNOR_STAGE_14 STAGE_13_OUT STAGE_14_INTERNAL STAGE_14_OUT VDD VDD GND GND NOR2_X1

XINV_STAGE_15 STAGE_16_OUT STAGE_15_INTERNAL VDD VDD GND GND INV_X1
XNOR_STAGE_15 STAGE_14_OUT STAGE_15_INTERNAL STAGE_15_OUT VDD VDD GND GND NOR2_X1

XINV_STAGE_16 STAGE_17_OUT STAGE_16_INTERNAL VDD VDD GND GND INV_X1
XNOR_STAGE_16 STAGE_15_OUT STAGE_16_INTERNAL STAGE_16_OUT VDD VDD GND GND NOR2_X1

XINV_STAGE_17 STAGE_18_OUT STAGE_17_INTERNAL VDD VDD GND GND INV_X1
XNOR_STAGE_17 STAGE_16_OUT STAGE_17_INTERNAL STAGE_17_OUT VDD VDD GND GND NOR2_X1

XINV_STAGE_18 STAGE_19_OUT STAGE_18_INTERNAL VDD VDD GND GND INV_X1
XNOR_STAGE_18 STAGE_17_OUT STAGE_18_INTERNAL STAGE_18_OUT VDD VDD GND GND NOR2_X1

XINV_STAGE_19 STAGE_20_OUT STAGE_19_INTERNAL VDD VDD GND GND INV_X1
XNOR_STAGE_19 STAGE_18_OUT STAGE_19_INTERNAL STAGE_19_OUT VDD VDD GND GND NOR2_X1

XINV_STAGE_20 STAGE_21_OUT STAGE_20_INTERNAL VDD VDD GND GND INV_X1
XNOR_STAGE_20 STAGE_19_OUT STAGE_20_INTERNAL STAGE_20_OUT VDD VDD GND GND NOR2_X1

XINV_STAGE_21 STAGE_22_OUT STAGE_21_INTERNAL VDD VDD GND GND INV_X1
XNOR_STAGE_21 STAGE_20_OUT STAGE_21_INTERNAL STAGE_21_OUT VDD VDD GND GND NOR2_X1

XINV_STAGE_22 STAGE_23_OUT STAGE_22_INTERNAL VDD VDD GND GND INV_X1
XNOR_STAGE_22 STAGE_21_OUT STAGE_22_INTERNAL STAGE_22_OUT VDD VDD GND GND NOR2_X1

XINV_STAGE_23 STAGE_24_OUT STAGE_23_INTERNAL VDD VDD GND GND INV_X1
XNOR_STAGE_23 STAGE_22_OUT STAGE_23_INTERNAL STAGE_23_OUT VDD VDD GND GND NOR2_X1

XINV_STAGE_24 STAGE_25_OUT STAGE_24_INTERNAL VDD VDD GND GND INV_X1
XNOR_STAGE_24 STAGE_23_OUT STAGE_24_INTERNAL STAGE_24_OUT VDD VDD GND GND NOR2_X1

XINV_STAGE_25 STAGE_26_OUT STAGE_25_INTERNAL VDD VDD GND GND INV_X1
XNOR_STAGE_25 STAGE_24_OUT STAGE_25_INTERNAL STAGE_25_OUT VDD VDD GND GND NOR2_X1

XINV_STAGE_26 STAGE_27_OUT STAGE_26_INTERNAL VDD VDD GND GND INV_X1
XNOR_STAGE_26 STAGE_25_OUT STAGE_26_INTERNAL STAGE_26_OUT VDD VDD GND GND NOR2_X1

XINV_STAGE_27 STAGE_28_OUT STAGE_27_INTERNAL VDD VDD GND GND INV_X1
XNOR_STAGE_27 STAGE_26_OUT STAGE_27_INTERNAL STAGE_27_OUT VDD VDD GND GND NOR2_X1

XINV_STAGE_28 STAGE_29_OUT STAGE_28_INTERNAL VDD VDD GND GND INV_X1
XNOR_STAGE_28 STAGE_27_OUT STAGE_28_INTERNAL STAGE_28_OUT VDD VDD GND GND NOR2_X1

XINV_STAGE_29 STAGE_0_OUT STAGE_29_INTERNAL VDD VDD GND GND INV_X1
XNOR_STAGE_29 STAGE_28_OUT STAGE_29_INTERNAL STAGE_29_OUT VDD VDD GND GND NOR2_X1


.PROBE TRAN V(PS_0_4)
.TRAN 0.1ps tend
.END
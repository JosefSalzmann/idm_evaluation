* circuit: nor inv chain
simulator lang=spice

.PARAM pw1=50ps pw2=400ps vsrc=0.8V srcdc=0.0V
*.PARAM pw1=50ps pw2=<sed>pw<sed>fs vsrc=supp srcdc=0.0V
.PARAM supp=0.8V slope=0.1fs start='0.1ns+pw1' realpw2='pw2-slope'
.PARAM t00=0.1ns t01='t00+0.2ns' t1='t01+0.4ns' t2='t1+6000fs' t3='t2+9000fs' t4='t3+8000fs'
.PARAM t5='t3+100000fs' t6='t5+100000fs'
.PARAM baseVal=0V peakVal=0.8V tend=2ns
*.PARAM baseVal=<sed>base<sed> peakVal=<sed>peak<sed>


.LIB /home/s11777724/involution_tool_library_files/backend/spice/fet.inc CMG

* main circuit
.INCLUDE /home/s11777724/involution_tool_library_files/backend/spice/cell/NOR2_X1.sp

**** SPECTRE Back Annotation
.option spef='../place_and_route/generic_parasitics.spef'
****

.TEMP 25
.OPTION
+ INGOLD=2
+ PARHIER=LOCAL
*+ POST=CSDF
+ PROBE
+ BRIEF
+ ACCURATE
+ ABSVAR=0.0001
+ DVDT=2
+ RELTOL=1e-11
*+ DELMAX=100fs
+ dc_pivot_check=yes

* vdd
VDD VDD GND 0.8v

VIN myin GND PWL 0ns baseVal t00 baseVal 't00+slope' peakVal t01 peakVal 't01+slope' baseVal 
+ t1 baseVal 't1+slope' peakVal t2 peakVal 't2+slope' baseVal
+ t3 baseVal 't3+slope' peakVal t4 peakVal 't4+slope' baseVal tend baseVal

XNOR0_1 myin GND STAGE0_1 VDD VDD GND GND NOR2_X1
* circuit under test
XNOR1_1 STAGE0_1 GND STAGE1_1 VDD VDD GND GND NOR2_X1
XNOR2_1 STAGE1_1 GND STAGE2_1 VDD VDD GND GND NOR2_X1
XNOR3_1 STAGE2_1 GND STAGE3_1 VDD VDD GND GND NOR2_X1
XNOR4_1 STAGE3_1 GND STAGE4_1 VDD VDD GND GND NOR2_X1
XNOR5_1 STAGE4_1 GND FANOUTTEST_1 VDD VDD GND GND NOR2_X1

XNOR5_1_1_1 FANOUTTEST_1 GND STAGE1_1_1 VDD VDD GND GND NOR2_X1
XNOR5_1_2_1 STAGE1_1_1 GND STAGE1_2_1 VDD VDD GND GND NOR2_X1
XNOR5_1_3_1 STAGE1_2_1 GND STAGE1_3_1 VDD VDD GND GND NOR2_X1
XNOR5_1_4_1 STAGE1_3_1 GND O_C_TERM1_4_1 VDD VDD GND GND NOR2_X1
C_TERM1_4_1 O_C_TERM1_4_1 GND 0.0779pF

XNOR5_2_1_1 FANOUTTEST_1 GND STAGE2_1_1 VDD VDD GND GND NOR2_X1
XNOR5_2_2_1 STAGE2_1_1 GND STAGE2_2_1 VDD VDD GND GND NOR2_X1
XNOR5_2_3_1 STAGE2_2_1 GND STAGE2_3_1 VDD VDD GND GND NOR2_X1
XNOR5_2_4_1 STAGE2_3_1 GND O_C_TERM2_4_1 VDD VDD GND GND NOR2_X1
C_TERM2_4_1 O_C_TERM2_4_1 GND 0.0779pF

XNOR5_3_1_1 FANOUTTEST_1 GND STAGE3_1_1 VDD VDD GND GND NOR2_X1
XNOR5_3_2_1 STAGE3_1_1 GND STAGE3_2_1 VDD VDD GND GND NOR2_X1
XNOR5_3_3_1 STAGE3_2_1 GND STAGE3_3_1 VDD VDD GND GND NOR2_X1
XNOR5_3_4_1 STAGE3_3_1 GND O_C_TERM3_4_1 VDD VDD GND GND NOR2_X1
C_TERM3_4_1 O_C_TERM3_4_1 GND 0.0779pF

XNOR5_4_1_1 FANOUTTEST_1 GND STAGE4_1_1 VDD VDD GND GND NOR2_X1
XNOR5_4_2_1 STAGE4_1_1 GND STAGE4_2_1 VDD VDD GND GND NOR2_X1
XNOR5_4_3_1 STAGE4_2_1 GND STAGE4_3_1 VDD VDD GND GND NOR2_X1
XNOR5_4_4_1 STAGE4_3_1 GND O_C_TERM4_4_1 VDD VDD GND GND NOR2_X1
C_TERM4_4_1 O_C_TERM4_4_1 GND 0.0779pF






XNOR0_2 myin GND STAGE0_2 VDD VDD GND GND NOR2_X1
XNOR1_2 STAGE0_2 GND STAGE1_2 VDD VDD GND GND NOR2_X1
XNOR2_2 STAGE1_2 GND STAGE2_2 VDD VDD GND GND NOR2_X1
XNOR3_2 STAGE2_2 GND STAGE3_2 VDD VDD GND GND NOR2_X1
XNOR4_2 STAGE3_2 GND STAGE4_2 VDD VDD GND GND NOR2_X1
XNOR5_2 STAGE4_2 GND FANOUTTEST_2 VDD VDD GND GND NOR2_X1

XNOR5_1_1_2 FANOUTTEST_2 VDD STAGE1_1_2 VDD VDD GND GND NOR2_X1
XNOR5_1_2_2 STAGE1_1_2 GND STAGE1_2_2 VDD VDD GND GND NOR2_X1
XNOR5_1_3_2 STAGE1_2_2 GND STAGE1_3_2 VDD VDD GND GND NOR2_X1
XNOR5_1_4_2 STAGE1_3_2 GND O_C_TERM1_4_2 VDD VDD GND GND NOR2_X1
C_TERM1_4_2 O_C_TERM1_4_2 GND 0.0779pF

XNOR5_2_1_2 FANOUTTEST_2 VDD STAGE2_1_2 VDD VDD GND GND NOR2_X1
XNOR5_2_2_2 STAGE2_1_2 GND STAGE2_2_2 VDD VDD GND GND NOR2_X1
XNOR5_2_3_2 STAGE2_2_2 GND STAGE2_3_2 VDD VDD GND GND NOR2_X1
XNOR5_2_4_2 STAGE2_3_2 GND O_C_TERM2_4_2 VDD VDD GND GND NOR2_X1
C_TERM2_4_2 O_C_TERM2_4_2 GND 0.0779pF

XNOR5_3_1_2 FANOUTTEST_2 GND STAGE3_1_2 VDD VDD GND GND NOR2_X1
XNOR5_3_2_2 STAGE3_1_2 GND STAGE3_2_2 VDD VDD GND GND NOR2_X1
XNOR5_3_3_2 STAGE3_2_2 GND STAGE3_3_2 VDD VDD GND GND NOR2_X1
XNOR5_3_4_2 STAGE3_3_2 GND O_C_TERM3_4_2 VDD VDD GND GND NOR2_X1
C_TERM3_4_2 O_C_TERM3_4_2 GND 0.0779pF

XNOR5_4_1_2 FANOUTTEST_2 GND STAGE4_1_2 VDD VDD GND GND NOR2_X1
XNOR5_4_2_2 STAGE4_1_2 GND STAGE4_2_2 VDD VDD GND GND NOR2_X1
XNOR5_4_3_2 STAGE4_2_2 GND STAGE4_3_2 VDD VDD GND GND NOR2_X1
XNOR5_4_4_2 STAGE4_3_2 GND O_C_TERM4_4_2 VDD VDD GND GND NOR2_X1
C_TERM4_4_2 O_C_TERM4_4_2 GND 0.0779pF





XNOR0_3 myin GND STAGE0_3 VDD VDD GND GND NOR2_X1
XNOR1_3 STAGE0_3 GND STAGE1_3 VDD VDD GND GND NOR2_X1
XNOR2_3 STAGE1_3 GND STAGE2_3 VDD VDD GND GND NOR2_X1
XNOR3_3 STAGE2_3 GND STAGE3_3 VDD VDD GND GND NOR2_X1
XNOR4_3 STAGE3_3 GND STAGE4_3 VDD VDD GND GND NOR2_X1
XNOR5_3 STAGE4_3 GND FANOUTTEST_3 VDD VDD GND GND NOR2_X1

XNOR5_1_1_3 FANOUTTEST_3 VDD STAGE1_1_3 VDD VDD GND GND NOR2_X1
XNOR5_1_2_3 STAGE1_1_3 GND STAGE1_2_3 VDD VDD GND GND NOR2_X1
XNOR5_1_3_3 STAGE1_2_3 GND STAGE1_3_3 VDD VDD GND GND NOR2_X1
XNOR5_1_4_3 STAGE1_3_3 GND O_C_TERM1_4_3 VDD VDD GND GND NOR2_X1
C_TERM1_4_3 O_C_TERM1_4_3 GND 0.0779pF

XNOR5_2_1_3 FANOUTTEST_3 VDD STAGE2_1_3 VDD VDD GND GND NOR2_X1
XNOR5_2_2_3 STAGE2_1_3 GND STAGE2_2_3 VDD VDD GND GND NOR2_X1
XNOR5_2_3_3 STAGE2_2_3 GND STAGE2_3_3 VDD VDD GND GND NOR2_X1
XNOR5_2_4_3 STAGE2_3_3 GND O_C_TERM2_4_3 VDD VDD GND GND NOR2_X1
C_TERM2_4_3 O_C_TERM2_4_3 GND 0.0779pF

XNOR5_3_1_3 FANOUTTEST_3 VDD STAGE3_1_3 VDD VDD GND GND NOR2_X1
XNOR5_3_2_3 STAGE3_1_3 GND STAGE3_2_3 VDD VDD GND GND NOR2_X1
XNOR5_3_3_3 STAGE3_2_3 GND STAGE3_3_3 VDD VDD GND GND NOR2_X1
XNOR5_3_4_3 STAGE3_3_3 GND O_C_TERM3_4_3 VDD VDD GND GND NOR2_X1
C_TERM3_4_3 O_C_TERM3_4_3 GND 0.0779pF

XNOR5_4_1_3 FANOUTTEST_3 VDD STAGE4_1_3 VDD VDD GND GND NOR2_X1
XNOR5_4_2_3 STAGE4_1_3 GND STAGE4_2_3 VDD VDD GND GND NOR2_X1
XNOR5_4_3_3 STAGE4_2_3 GND STAGE4_3_3 VDD VDD GND GND NOR2_X1
XNOR5_4_4_3 STAGE4_3_3 GND O_C_TERM4_4_3 VDD VDD GND GND NOR2_X1
C_TERM4_4_3 O_C_TERM4_4_3 GND 0.0779pF





.PROBE TRAN V(myin) V(STAGE4_1) V(STAGE4_2) V(STAGE4_3) V(FANOUTTEST_1) V(FANOUTTEST_2) V(FANOUTTEST_3)
.TRAN 0.1ps tend
.END

module nor_inv_chain_100_stages (myin, myout);
       input myin;
       output myout;

       wire GND = 1'b0;
       wire STAGE0, STAGE1, STAGE2, STAGE3, STAGE4, STAGE5, STAGE6, STAGE7, STAGE8, STAGE9, STAGE10, STAGE11, STAGE12, STAGE13, STAGE14, STAGE15, STAGE16, STAGE17, STAGE18, STAGE19, STAGE20, STAGE21, STAGE22, STAGE23, STAGE24, STAGE25, STAGE26, STAGE27, STAGE28, STAGE29, STAGE30, STAGE31, STAGE32, STAGE33, STAGE34, STAGE35, STAGE36, STAGE37, STAGE38, STAGE39, STAGE40, STAGE41, STAGE42, STAGE43, STAGE44, STAGE45, STAGE46, STAGE47, STAGE48, STAGE49, STAGE50, STAGE51, STAGE52, STAGE53, STAGE54, STAGE55, STAGE56, STAGE57, STAGE58, STAGE59, STAGE60, STAGE61, STAGE62, STAGE63, STAGE64, STAGE65, STAGE66, STAGE67, STAGE68, STAGE69, STAGE70, STAGE71, STAGE72, STAGE73, STAGE74, STAGE75, STAGE76, STAGE77, STAGE78, STAGE79, STAGE80, STAGE81, STAGE82, STAGE83, STAGE84, STAGE85, STAGE86, STAGE87, STAGE88, STAGE89, STAGE90, STAGE91, STAGE92, STAGE93, STAGE94, STAGE95, STAGE96, STAGE97, STAGE98, STAGE99, STAGE100, STAGE101, STAGE102, STAGE103, STAGE104, STAGE105, STAGE106, STAGE107, STAGE108, STAGE109, STAGE110, STAGE111, STAGE112, STAGE113, STAGE114, STAGE115, STAGE116, STAGE117, STAGE118, STAGE119;


       NOR2_X1 NOR0 ( .A1 (myin), .A2 (GND), .ZN (STAGE0));
       NOR2_X1 NOR1 ( .A1 (STAGE0), .A2 (GND), .ZN (STAGE1));   
       NOR2_X1 NOR2 ( .A1 (STAGE1), .A2 (GND), .ZN (STAGE2));   
       NOR2_X1 NOR3 ( .A1 (STAGE2), .A2 (GND), .ZN (STAGE3));   
       NOR2_X1 NOR4 ( .A1 (STAGE3), .A2 (GND), .ZN (STAGE4));   
       NOR2_X1 NOR5 ( .A1 (STAGE4), .A2 (GND), .ZN (STAGE5));   
       NOR2_X1 NOR6 ( .A1 (STAGE5), .A2 (GND), .ZN (STAGE6));   
       NOR2_X1 NOR7 ( .A1 (STAGE6), .A2 (GND), .ZN (STAGE7));   
       NOR2_X1 NOR8 ( .A1 (STAGE7), .A2 (GND), .ZN (STAGE8));   
       NOR2_X1 NOR9 ( .A1 (STAGE8), .A2 (GND), .ZN (STAGE9));   
       NOR2_X1 NOR10 ( .A1 (STAGE9), .A2 (GND), .ZN (STAGE10)); 
       NOR2_X1 NOR11 ( .A1 (STAGE10), .A2 (GND), .ZN (STAGE11));
       NOR2_X1 NOR12 ( .A1 (STAGE11), .A2 (GND), .ZN (STAGE12));
       NOR2_X1 NOR13 ( .A1 (STAGE12), .A2 (GND), .ZN (STAGE13));
       NOR2_X1 NOR14 ( .A1 (STAGE13), .A2 (GND), .ZN (STAGE14));
       NOR2_X1 NOR15 ( .A1 (STAGE14), .A2 (GND), .ZN (STAGE15));
       NOR2_X1 NOR16 ( .A1 (STAGE15), .A2 (GND), .ZN (STAGE16));
       NOR2_X1 NOR17 ( .A1 (STAGE16), .A2 (GND), .ZN (STAGE17));
       NOR2_X1 NOR18 ( .A1 (STAGE17), .A2 (GND), .ZN (STAGE18));
       NOR2_X1 NOR19 ( .A1 (STAGE18), .A2 (GND), .ZN (STAGE19));
       NOR2_X1 NOR20 ( .A1 (STAGE19), .A2 (GND), .ZN (STAGE20));
       NOR2_X1 NOR21 ( .A1 (STAGE20), .A2 (GND), .ZN (STAGE21));
       NOR2_X1 NOR22 ( .A1 (STAGE21), .A2 (GND), .ZN (STAGE22));
       NOR2_X1 NOR23 ( .A1 (STAGE22), .A2 (GND), .ZN (STAGE23));
       NOR2_X1 NOR24 ( .A1 (STAGE23), .A2 (GND), .ZN (STAGE24));
       NOR2_X1 NOR25 ( .A1 (STAGE24), .A2 (GND), .ZN (STAGE25));
       NOR2_X1 NOR26 ( .A1 (STAGE25), .A2 (GND), .ZN (STAGE26));
       NOR2_X1 NOR27 ( .A1 (STAGE26), .A2 (GND), .ZN (STAGE27));
       NOR2_X1 NOR28 ( .A1 (STAGE27), .A2 (GND), .ZN (STAGE28));
       NOR2_X1 NOR29 ( .A1 (STAGE28), .A2 (GND), .ZN (STAGE29));
       NOR2_X1 NOR30 ( .A1 (STAGE29), .A2 (GND), .ZN (STAGE30));
       NOR2_X1 NOR31 ( .A1 (STAGE30), .A2 (GND), .ZN (STAGE31));
       NOR2_X1 NOR32 ( .A1 (STAGE31), .A2 (GND), .ZN (STAGE32));
       NOR2_X1 NOR33 ( .A1 (STAGE32), .A2 (GND), .ZN (STAGE33));
       NOR2_X1 NOR34 ( .A1 (STAGE33), .A2 (GND), .ZN (STAGE34));
       NOR2_X1 NOR35 ( .A1 (STAGE34), .A2 (GND), .ZN (STAGE35));
       NOR2_X1 NOR36 ( .A1 (STAGE35), .A2 (GND), .ZN (STAGE36));
       NOR2_X1 NOR37 ( .A1 (STAGE36), .A2 (GND), .ZN (STAGE37));
       NOR2_X1 NOR38 ( .A1 (STAGE37), .A2 (GND), .ZN (STAGE38));
       NOR2_X1 NOR39 ( .A1 (STAGE38), .A2 (GND), .ZN (STAGE39));
       NOR2_X1 NOR40 ( .A1 (STAGE39), .A2 (GND), .ZN (STAGE40));
       NOR2_X1 NOR41 ( .A1 (STAGE40), .A2 (GND), .ZN (STAGE41));
       NOR2_X1 NOR42 ( .A1 (STAGE41), .A2 (GND), .ZN (STAGE42));
       NOR2_X1 NOR43 ( .A1 (STAGE42), .A2 (GND), .ZN (STAGE43));
       NOR2_X1 NOR44 ( .A1 (STAGE43), .A2 (GND), .ZN (STAGE44));
       NOR2_X1 NOR45 ( .A1 (STAGE44), .A2 (GND), .ZN (STAGE45));
       NOR2_X1 NOR46 ( .A1 (STAGE45), .A2 (GND), .ZN (STAGE46));
       NOR2_X1 NOR47 ( .A1 (STAGE46), .A2 (GND), .ZN (STAGE47));
       NOR2_X1 NOR48 ( .A1 (STAGE47), .A2 (GND), .ZN (STAGE48));
       NOR2_X1 NOR49 ( .A1 (STAGE48), .A2 (GND), .ZN (STAGE49));
       NOR2_X1 NOR50 ( .A1 (STAGE49), .A2 (GND), .ZN (STAGE50));
       NOR2_X1 NOR51 ( .A1 (STAGE50), .A2 (GND), .ZN (STAGE51));
       NOR2_X1 NOR52 ( .A1 (STAGE51), .A2 (GND), .ZN (STAGE52));
       NOR2_X1 NOR53 ( .A1 (STAGE52), .A2 (GND), .ZN (STAGE53));
       NOR2_X1 NOR54 ( .A1 (STAGE53), .A2 (GND), .ZN (STAGE54));
       NOR2_X1 NOR55 ( .A1 (STAGE54), .A2 (GND), .ZN (STAGE55));
       NOR2_X1 NOR56 ( .A1 (STAGE55), .A2 (GND), .ZN (STAGE56));
       NOR2_X1 NOR57 ( .A1 (STAGE56), .A2 (GND), .ZN (STAGE57));
       NOR2_X1 NOR58 ( .A1 (STAGE57), .A2 (GND), .ZN (STAGE58));
       NOR2_X1 NOR59 ( .A1 (STAGE58), .A2 (GND), .ZN (STAGE59));
       NOR2_X1 NOR60 ( .A1 (STAGE59), .A2 (GND), .ZN (STAGE60));
       NOR2_X1 NOR61 ( .A1 (STAGE60), .A2 (GND), .ZN (STAGE61));
       NOR2_X1 NOR62 ( .A1 (STAGE61), .A2 (GND), .ZN (STAGE62));
       NOR2_X1 NOR63 ( .A1 (STAGE62), .A2 (GND), .ZN (STAGE63));
       NOR2_X1 NOR64 ( .A1 (STAGE63), .A2 (GND), .ZN (STAGE64));
       NOR2_X1 NOR65 ( .A1 (STAGE64), .A2 (GND), .ZN (STAGE65));
       NOR2_X1 NOR66 ( .A1 (STAGE65), .A2 (GND), .ZN (STAGE66));
       NOR2_X1 NOR67 ( .A1 (STAGE66), .A2 (GND), .ZN (STAGE67));
       NOR2_X1 NOR68 ( .A1 (STAGE67), .A2 (GND), .ZN (STAGE68));
       NOR2_X1 NOR69 ( .A1 (STAGE68), .A2 (GND), .ZN (STAGE69));
       NOR2_X1 NOR70 ( .A1 (STAGE69), .A2 (GND), .ZN (STAGE70));
       NOR2_X1 NOR71 ( .A1 (STAGE70), .A2 (GND), .ZN (STAGE71));
       NOR2_X1 NOR72 ( .A1 (STAGE71), .A2 (GND), .ZN (STAGE72));
       NOR2_X1 NOR73 ( .A1 (STAGE72), .A2 (GND), .ZN (STAGE73));
       NOR2_X1 NOR74 ( .A1 (STAGE73), .A2 (GND), .ZN (STAGE74));
       NOR2_X1 NOR75 ( .A1 (STAGE74), .A2 (GND), .ZN (STAGE75));
       NOR2_X1 NOR76 ( .A1 (STAGE75), .A2 (GND), .ZN (STAGE76));
       NOR2_X1 NOR77 ( .A1 (STAGE76), .A2 (GND), .ZN (STAGE77));
       NOR2_X1 NOR78 ( .A1 (STAGE77), .A2 (GND), .ZN (STAGE78));
       NOR2_X1 NOR79 ( .A1 (STAGE78), .A2 (GND), .ZN (STAGE79));
       NOR2_X1 NOR80 ( .A1 (STAGE79), .A2 (GND), .ZN (STAGE80));
       NOR2_X1 NOR81 ( .A1 (STAGE80), .A2 (GND), .ZN (STAGE81));
       NOR2_X1 NOR82 ( .A1 (STAGE81), .A2 (GND), .ZN (STAGE82));
       NOR2_X1 NOR83 ( .A1 (STAGE82), .A2 (GND), .ZN (STAGE83));
       NOR2_X1 NOR84 ( .A1 (STAGE83), .A2 (GND), .ZN (STAGE84));
       NOR2_X1 NOR85 ( .A1 (STAGE84), .A2 (GND), .ZN (STAGE85));
       NOR2_X1 NOR86 ( .A1 (STAGE85), .A2 (GND), .ZN (STAGE86));
       NOR2_X1 NOR87 ( .A1 (STAGE86), .A2 (GND), .ZN (STAGE87));
       NOR2_X1 NOR88 ( .A1 (STAGE87), .A2 (GND), .ZN (STAGE88));
       NOR2_X1 NOR89 ( .A1 (STAGE88), .A2 (GND), .ZN (STAGE89));
       NOR2_X1 NOR90 ( .A1 (STAGE89), .A2 (GND), .ZN (STAGE90));
       NOR2_X1 NOR91 ( .A1 (STAGE90), .A2 (GND), .ZN (STAGE91));
       NOR2_X1 NOR92 ( .A1 (STAGE91), .A2 (GND), .ZN (STAGE92));
       NOR2_X1 NOR93 ( .A1 (STAGE92), .A2 (GND), .ZN (STAGE93));
       NOR2_X1 NOR94 ( .A1 (STAGE93), .A2 (GND), .ZN (STAGE94));
       NOR2_X1 NOR95 ( .A1 (STAGE94), .A2 (GND), .ZN (STAGE95));
       NOR2_X1 NOR96 ( .A1 (STAGE95), .A2 (GND), .ZN (STAGE96));
       NOR2_X1 NOR97 ( .A1 (STAGE96), .A2 (GND), .ZN (STAGE97));
       NOR2_X1 NOR98 ( .A1 (STAGE97), .A2 (GND), .ZN (STAGE98));
       NOR2_X1 NOR99 ( .A1 (STAGE98), .A2 (GND), .ZN (STAGE99));
       NOR2_X1 NOR100 ( .A1 (STAGE99), .A2 (GND), .ZN (STAGE100));
       NOR2_X1 NOR101 ( .A1 (STAGE100), .A2 (GND), .ZN (STAGE101));
       NOR2_X1 NOR102 ( .A1 (STAGE101), .A2 (GND), .ZN (STAGE102));
       NOR2_X1 NOR103 ( .A1 (STAGE102), .A2 (GND), .ZN (STAGE103));
       NOR2_X1 NOR104 ( .A1 (STAGE103), .A2 (GND), .ZN (STAGE104));
       NOR2_X1 NOR105 ( .A1 (STAGE104), .A2 (GND), .ZN (STAGE105));
       NOR2_X1 NOR106 ( .A1 (STAGE105), .A2 (GND), .ZN (STAGE106));
       NOR2_X1 NOR107 ( .A1 (STAGE106), .A2 (GND), .ZN (STAGE107));
       NOR2_X1 NOR108 ( .A1 (STAGE107), .A2 (GND), .ZN (STAGE108));
       NOR2_X1 NOR109 ( .A1 (STAGE108), .A2 (GND), .ZN (STAGE109));
       NOR2_X1 NOR110 ( .A1 (STAGE109), .A2 (GND), .ZN (STAGE110));
       NOR2_X1 NOR111 ( .A1 (STAGE110), .A2 (GND), .ZN (STAGE111));
       NOR2_X1 NOR112 ( .A1 (STAGE111), .A2 (GND), .ZN (STAGE112));
       NOR2_X1 NOR113 ( .A1 (STAGE112), .A2 (GND), .ZN (STAGE113));
       NOR2_X1 NOR114 ( .A1 (STAGE113), .A2 (GND), .ZN (STAGE114));
       NOR2_X1 NOR115 ( .A1 (STAGE114), .A2 (GND), .ZN (STAGE115));
       NOR2_X1 NOR116 ( .A1 (STAGE115), .A2 (GND), .ZN (STAGE116));
       NOR2_X1 NOR117 ( .A1 (STAGE116), .A2 (GND), .ZN (STAGE117));
       NOR2_X1 NOR118 ( .A1 (STAGE117), .A2 (GND), .ZN (STAGE118));
       NOR2_X1 NOR119 ( .A1 (STAGE118), .A2 (GND), .ZN (myout));

endmodule

module c17_NOR_template (N1_PWL, N2_PWL, N3_PWL, N6_PWL, N7_PWL, N22_TERMINATION, N23_TERMINATION);
       input N1_PWL, N2_PWL, N3_PWL, N6_PWL, N7_PWL;
       output N22_TERMINATION, N23_TERMINATION;

       wire GND = 1'b0;
       wire XNOR_1_1_N1_PULSESHAPING_OUT, XNOR_1_2_N1_PULSESHAPING_OUT, XNOR_1_3_N1_PULSESHAPING_OUT, XNOR_1_4_N1_PULSESHAPING_OUT, XNOR_1_5_N1_PULSESHAPING_OUT, XNOR_1_6_N1_PULSESHAPING_OUT;
       NOR2_X1 XNOR_1_1_N1_PULSESHAPING (.ZN (XNOR_1_1_N1_PULSESHAPING_OUT), .A1 (N1_PWL), .A2 (GND));
       NOR2_X1 XNOR_1_2_N1_PULSESHAPING (.ZN (XNOR_1_2_N1_PULSESHAPING_OUT), .A1 (XNOR_1_1_N1_PULSESHAPING_OUT), .A2 (GND));
       NOR2_X1 XNOR_1_3_N1_PULSESHAPING (.ZN (XNOR_1_3_N1_PULSESHAPING_OUT), .A1 (XNOR_1_2_N1_PULSESHAPING_OUT), .A2 (GND));
       NOR2_X1 XNOR_1_4_N1_PULSESHAPING (.ZN (XNOR_1_4_N1_PULSESHAPING_OUT), .A1 (XNOR_1_3_N1_PULSESHAPING_OUT), .A2 (GND));
       NOR2_X1 XNOR_1_5_N1_PULSESHAPING (.ZN (XNOR_1_5_N1_PULSESHAPING_OUT), .A1 (XNOR_1_4_N1_PULSESHAPING_OUT), .A2 (GND));
       NOR2_X1 XNOR_1_6_N1_PULSESHAPING (.ZN (XNOR_1_6_N1_PULSESHAPING_OUT), .A1 (XNOR_1_5_N1_PULSESHAPING_OUT), .A2 (GND));
       NOR2_X1 XNOR_1_7_N1_PULSESHAPING (.ZN (N1), .A1 (XNOR_1_6_N1_PULSESHAPING_OUT), .A2 (GND));

       wire XNOR_1_1_N2_PULSESHAPING_OUT, XNOR_1_2_N2_PULSESHAPING_OUT, XNOR_1_3_N2_PULSESHAPING_OUT, XNOR_1_4_N2_PULSESHAPING_OUT, XNOR_1_5_N2_PULSESHAPING_OUT, XNOR_1_6_N2_PULSESHAPING_OUT;
       NOR2_X1 XNOR_1_1_N2_PULSESHAPING (.ZN (XNOR_1_1_N2_PULSESHAPING_OUT), .A1 (N2_PWL), .A2 (GND));
       NOR2_X1 XNOR_1_2_N2_PULSESHAPING (.ZN (XNOR_1_2_N2_PULSESHAPING_OUT), .A1 (XNOR_1_1_N2_PULSESHAPING_OUT), .A2 (GND));
       NOR2_X1 XNOR_1_3_N2_PULSESHAPING (.ZN (XNOR_1_3_N2_PULSESHAPING_OUT), .A1 (XNOR_1_2_N2_PULSESHAPING_OUT), .A2 (GND));
       NOR2_X1 XNOR_1_4_N2_PULSESHAPING (.ZN (XNOR_1_4_N2_PULSESHAPING_OUT), .A1 (XNOR_1_3_N2_PULSESHAPING_OUT), .A2 (GND));
       NOR2_X1 XNOR_1_5_N2_PULSESHAPING (.ZN (XNOR_1_5_N2_PULSESHAPING_OUT), .A1 (XNOR_1_4_N2_PULSESHAPING_OUT), .A2 (GND));
       NOR2_X1 XNOR_1_6_N2_PULSESHAPING (.ZN (XNOR_1_6_N2_PULSESHAPING_OUT), .A1 (XNOR_1_5_N2_PULSESHAPING_OUT), .A2 (GND));
       NOR2_X1 XNOR_1_7_N2_PULSESHAPING (.ZN (N2), .A1 (XNOR_1_6_N2_PULSESHAPING_OUT), .A2 (GND));

       wire XNOR_1_1_N3_PULSESHAPING_OUT, XNOR_1_2_N3_PULSESHAPING_OUT, XNOR_1_3_N3_PULSESHAPING_OUT, XNOR_1_4_N3_PULSESHAPING_OUT, XNOR_1_5_N3_PULSESHAPING_OUT, XNOR_1_6_N3_PULSESHAPING_OUT;
       NOR2_X1 XNOR_1_1_N3_PULSESHAPING (.ZN (XNOR_1_1_N3_PULSESHAPING_OUT), .A1 (N3_PWL), .A2 (GND));
       NOR2_X1 XNOR_1_2_N3_PULSESHAPING (.ZN (XNOR_1_2_N3_PULSESHAPING_OUT), .A1 (XNOR_1_1_N3_PULSESHAPING_OUT), .A2 (GND));
       NOR2_X1 XNOR_1_3_N3_PULSESHAPING (.ZN (XNOR_1_3_N3_PULSESHAPING_OUT), .A1 (XNOR_1_2_N3_PULSESHAPING_OUT), .A2 (GND));
       NOR2_X1 XNOR_1_4_N3_PULSESHAPING (.ZN (XNOR_1_4_N3_PULSESHAPING_OUT), .A1 (XNOR_1_3_N3_PULSESHAPING_OUT), .A2 (GND));
       NOR2_X1 XNOR_1_5_N3_PULSESHAPING (.ZN (XNOR_1_5_N3_PULSESHAPING_OUT), .A1 (XNOR_1_4_N3_PULSESHAPING_OUT), .A2 (GND));
       NOR2_X1 XNOR_1_6_N3_PULSESHAPING (.ZN (XNOR_1_6_N3_PULSESHAPING_OUT), .A1 (XNOR_1_5_N3_PULSESHAPING_OUT), .A2 (GND));
       NOR2_X1 XNOR_1_7_N3_PULSESHAPING (.ZN (N3), .A1 (XNOR_1_6_N3_PULSESHAPING_OUT), .A2 (GND));

       wire XNOR_1_1_N6_PULSESHAPING_OUT, XNOR_1_2_N6_PULSESHAPING_OUT, XNOR_1_3_N6_PULSESHAPING_OUT, XNOR_1_4_N6_PULSESHAPING_OUT, XNOR_1_5_N6_PULSESHAPING_OUT, XNOR_1_6_N6_PULSESHAPING_OUT;
       NOR2_X1 XNOR_1_1_N6_PULSESHAPING (.ZN (XNOR_1_1_N6_PULSESHAPING_OUT), .A1 (N6_PWL), .A2 (GND));
       NOR2_X1 XNOR_1_2_N6_PULSESHAPING (.ZN (XNOR_1_2_N6_PULSESHAPING_OUT), .A1 (XNOR_1_1_N6_PULSESHAPING_OUT), .A2 (GND));
       NOR2_X1 XNOR_1_3_N6_PULSESHAPING (.ZN (XNOR_1_3_N6_PULSESHAPING_OUT), .A1 (XNOR_1_2_N6_PULSESHAPING_OUT), .A2 (GND));
       NOR2_X1 XNOR_1_4_N6_PULSESHAPING (.ZN (XNOR_1_4_N6_PULSESHAPING_OUT), .A1 (XNOR_1_3_N6_PULSESHAPING_OUT), .A2 (GND));
       NOR2_X1 XNOR_1_5_N6_PULSESHAPING (.ZN (XNOR_1_5_N6_PULSESHAPING_OUT), .A1 (XNOR_1_4_N6_PULSESHAPING_OUT), .A2 (GND));
       NOR2_X1 XNOR_1_6_N6_PULSESHAPING (.ZN (XNOR_1_6_N6_PULSESHAPING_OUT), .A1 (XNOR_1_5_N6_PULSESHAPING_OUT), .A2 (GND));
       NOR2_X1 XNOR_1_7_N6_PULSESHAPING (.ZN (N6), .A1 (XNOR_1_6_N6_PULSESHAPING_OUT), .A2 (GND));

       wire XNOR_1_1_N7_PULSESHAPING_OUT, XNOR_1_2_N7_PULSESHAPING_OUT, XNOR_1_3_N7_PULSESHAPING_OUT, XNOR_1_4_N7_PULSESHAPING_OUT, XNOR_1_5_N7_PULSESHAPING_OUT, XNOR_1_6_N7_PULSESHAPING_OUT;
       NOR2_X1 XNOR_1_1_N7_PULSESHAPING (.ZN (XNOR_1_1_N7_PULSESHAPING_OUT), .A1 (N7_PWL), .A2 (GND));
       NOR2_X1 XNOR_1_2_N7_PULSESHAPING (.ZN (XNOR_1_2_N7_PULSESHAPING_OUT), .A1 (XNOR_1_1_N7_PULSESHAPING_OUT), .A2 (GND));
       NOR2_X1 XNOR_1_3_N7_PULSESHAPING (.ZN (XNOR_1_3_N7_PULSESHAPING_OUT), .A1 (XNOR_1_2_N7_PULSESHAPING_OUT), .A2 (GND));
       NOR2_X1 XNOR_1_4_N7_PULSESHAPING (.ZN (XNOR_1_4_N7_PULSESHAPING_OUT), .A1 (XNOR_1_3_N7_PULSESHAPING_OUT), .A2 (GND));
       NOR2_X1 XNOR_1_5_N7_PULSESHAPING (.ZN (XNOR_1_5_N7_PULSESHAPING_OUT), .A1 (XNOR_1_4_N7_PULSESHAPING_OUT), .A2 (GND));
       NOR2_X1 XNOR_1_6_N7_PULSESHAPING (.ZN (XNOR_1_6_N7_PULSESHAPING_OUT), .A1 (XNOR_1_5_N7_PULSESHAPING_OUT), .A2 (GND));
       NOR2_X1 XNOR_1_7_N7_PULSESHAPING (.ZN (N7), .A1 (XNOR_1_6_N7_PULSESHAPING_OUT), .A2 (GND));



       wire XNOR_1_1_NUM1_OUT, XNOR_1_2_NUM1_OUT, XNOR_1_3_NUM1_OUT;
       NOR2_X1 XNOR_1_1_NUM1 (.ZN (XNOR_1_1_NUM1_OUT), .A1 (N1), .A2 (GND));
       NOR2_X1 XNOR_1_2_NUM1 (.ZN (XNOR_1_2_NUM1_OUT), .A1 (GND), .A2 (N3));
       NOR2_X1 XNOR_1_3_NUM1 (.ZN (XNOR_1_3_NUM1_OUT), .A1 (XNOR_1_1_NUM1_OUT), .A2 (XNOR_1_2_NUM1_OUT));
       NOR2_X1 XNOR_1_4_NUM1 (.ZN (N10), .A1 (XNOR_1_3_NUM1_OUT), .A2 (GND));
       wire XNOR_1_1_NUM2_OUT, XNOR_1_2_NUM2_OUT, XNOR_1_3_NUM2_OUT;
       NOR2_X1 XNOR_1_1_NUM2 (.ZN (XNOR_1_1_NUM2_OUT), .A1 (N3), .A2 (GND));
       NOR2_X1 XNOR_1_2_NUM2 (.ZN (XNOR_1_2_NUM2_OUT), .A1 (GND), .A2 (N6));
       NOR2_X1 XNOR_1_3_NUM2 (.ZN (XNOR_1_3_NUM2_OUT), .A1 (XNOR_1_1_NUM2_OUT), .A2 (XNOR_1_2_NUM2_OUT));
       NOR2_X1 XNOR_1_4_NUM2 (.ZN (N11), .A1 (XNOR_1_3_NUM2_OUT), .A2 (GND));
       wire XNOR_1_1_NUM3_OUT, XNOR_1_2_NUM3_OUT, XNOR_1_3_NUM3_OUT;
       NOR2_X1 XNOR_1_1_NUM3 (.ZN (XNOR_1_1_NUM3_OUT), .A1 (N2), .A2 (GND));
       NOR2_X1 XNOR_1_2_NUM3 (.ZN (XNOR_1_2_NUM3_OUT), .A1 (GND), .A2 (N11));
       NOR2_X1 XNOR_1_3_NUM3 (.ZN (XNOR_1_3_NUM3_OUT), .A1 (XNOR_1_1_NUM3_OUT), .A2 (XNOR_1_2_NUM3_OUT));
       NOR2_X1 XNOR_1_4_NUM3 (.ZN (N16), .A1 (XNOR_1_3_NUM3_OUT), .A2 (GND));
       wire XNOR_1_1_NUM4_OUT, XNOR_1_2_NUM4_OUT, XNOR_1_3_NUM4_OUT;
       NOR2_X1 XNOR_1_1_NUM4 (.ZN (XNOR_1_1_NUM4_OUT), .A1 (N11), .A2 (GND));
       NOR2_X1 XNOR_1_2_NUM4 (.ZN (XNOR_1_2_NUM4_OUT), .A1 (GND), .A2 (N7));
       NOR2_X1 XNOR_1_3_NUM4 (.ZN (XNOR_1_3_NUM4_OUT), .A1 (XNOR_1_1_NUM4_OUT), .A2 (XNOR_1_2_NUM4_OUT));
       NOR2_X1 XNOR_1_4_NUM4 (.ZN (N19), .A1 (XNOR_1_3_NUM4_OUT), .A2 (GND));
       wire XNOR_1_1_NUM5_OUT, XNOR_1_2_NUM5_OUT, XNOR_1_3_NUM5_OUT;
       NOR2_X1 XNOR_1_1_NUM5 (.ZN (XNOR_1_1_NUM5_OUT), .A1 (N10), .A2 (GND));
       NOR2_X1 XNOR_1_2_NUM5 (.ZN (XNOR_1_2_NUM5_OUT), .A1 (GND), .A2 (N16));
       NOR2_X1 XNOR_1_3_NUM5 (.ZN (XNOR_1_3_NUM5_OUT), .A1 (XNOR_1_1_NUM5_OUT), .A2 (XNOR_1_2_NUM5_OUT));
       NOR2_X1 XNOR_1_4_NUM5 (.ZN (N22), .A1 (XNOR_1_3_NUM5_OUT), .A2 (GND));
       wire XNOR_1_1_NUM6_OUT, XNOR_1_2_NUM6_OUT, XNOR_1_3_NUM6_OUT;
       NOR2_X1 XNOR_1_1_NUM6 (.ZN (XNOR_1_1_NUM6_OUT), .A1 (N16), .A2 (GND));
       NOR2_X1 XNOR_1_2_NUM6 (.ZN (XNOR_1_2_NUM6_OUT), .A1 (GND), .A2 (N19));
       NOR2_X1 XNOR_1_3_NUM6 (.ZN (XNOR_1_3_NUM6_OUT), .A1 (XNOR_1_1_NUM6_OUT), .A2 (XNOR_1_2_NUM6_OUT));
       NOR2_X1 XNOR_1_4_NUM6 (.ZN (N23), .A1 (XNOR_1_3_NUM6_OUT), .A2 (GND));


       wire XNOR_1_1_N22_TERMINATION_OUT, XNOR_1_2_N22_TERMINATION_OUT;
       NOR2_X1 XNOR_1_1_N22_TERMINATION (.ZN (XNOR_1_1_N22_TERMINATION_OUT), .A1 (N22), .A2 (GND));
       NOR2_X1 XNOR_1_2_N22_TERMINATION (.ZN (N22_TERMINATION), .A1 (XNOR_1_1_N22_TERMINATION_OUT), .A2 (XNOR_1_2_N22_TERMINATION_OUT));

       wire XNOR_1_1_N23_TERMINATION_OUT, XNOR_1_2_N23_TERMINATION_OUT;
       NOR2_X1 XNOR_1_1_N23_TERMINATION (.ZN (XNOR_1_1_N23_TERMINATION_OUT), .A1 (N23), .A2 (GND));
       NOR2_X1 XNOR_1_2_N23_TERMINATION (.ZN (N23_TERMINATION), .A1 (XNOR_1_1_N23_TERMINATION_OUT), .A2 (XNOR_1_2_N23_TERMINATION_OUT));



endmodule
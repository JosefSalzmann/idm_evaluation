* circuit: nor inv chain
simulator lang=spice

*.PARAM pw=<sed>pw<sed>as
.PARAM supp=0.8V slope=0.1fs
.PARAM t_init0=0.1ns t_init1=0.174ns
.PARAM baseVal=0V peakVal=0.8V tend=1.0ns


.LIB /home/s11777724/involution_tool_library_files/backend/spice/fet.inc CMG

* main circuit
.INCLUDE /home/s11777724/involution_tool_library_files/backend/spice/cell/NOR2_X1.sp

**** SPECTRE Back Annotation
.option spef='../place_and_route/generic_parasitics.spef'
****

.TEMP 25
.OPTION
+ INGOLD=2
+ PARHIER=LOCAL
*+ POST=CSDF
+ PROBE
+ BRIEF
+ ACCURATE
+ ABSVAR=0.0001
+ DVDT=2
+ RELTOL=1e-11
*+ DELMAX=100fs
+ dc_pivot_check=yes

* vdd
VDD VDD GND 0.8v

VIN myin GND PWL 0ns baseVal t_init0 baseVal 't_init0+slope' peakVal t_init1 peakVal 't_init1+slope' baseVal

* circuit under test
XNOR0 myin GND STAGE0 VDD VDD GND GND NOR2_X1
XNOR1 STAGE0 GND STAGE1 VDD VDD GND GND NOR2_X1
XNOR2 STAGE1 GND STAGE2 VDD VDD GND GND NOR2_X1
XNOR3 STAGE2 GND STAGE3 VDD VDD GND GND NOR2_X1
XNOR4 STAGE3 GND STAGE4 VDD VDD GND GND NOR2_X1
XNOR5 STAGE4 GND STAGE5 VDD VDD GND GND NOR2_X1
XNOR6 STAGE5 GND STAGE6 VDD VDD GND GND NOR2_X1
XNOR7 STAGE6 GND STAGE7 VDD VDD GND GND NOR2_X1
XNOR8 STAGE7 GND STAGE8 VDD VDD GND GND NOR2_X1
XNOR9 STAGE8 GND STAGE9 VDD VDD GND GND NOR2_X1
XNOR10 STAGE9 GND STAGE10 VDD VDD GND GND NOR2_X1
XNOR11 STAGE10 GND STAGE11 VDD VDD GND GND NOR2_X1
XNOR12 STAGE11 GND STAGE12 VDD VDD GND GND NOR2_X1
XNOR13 STAGE12 GND STAGE13 VDD VDD GND GND NOR2_X1
XNOR14 STAGE13 GND STAGE14 VDD VDD GND GND NOR2_X1
XNOR15 STAGE14 GND STAGE15 VDD VDD GND GND NOR2_X1
XNOR16 STAGE15 GND STAGE16 VDD VDD GND GND NOR2_X1
XNOR17 STAGE16 GND STAGE17 VDD VDD GND GND NOR2_X1
XNOR18 STAGE17 GND STAGE18 VDD VDD GND GND NOR2_X1
XNOR19 STAGE18 GND STAGE19 VDD VDD GND GND NOR2_X1
XNOR20 STAGE19 GND STAGE20 VDD VDD GND GND NOR2_X1
XNOR21 STAGE20 GND STAGE21 VDD VDD GND GND NOR2_X1
XNOR22 STAGE21 GND STAGE22 VDD VDD GND GND NOR2_X1
XNOR23 STAGE22 GND STAGE23 VDD VDD GND GND NOR2_X1
XNOR24 STAGE23 GND STAGE24 VDD VDD GND GND NOR2_X1
XNOR25 STAGE24 GND STAGE25 VDD VDD GND GND NOR2_X1
XNOR26 STAGE25 GND STAGE26 VDD VDD GND GND NOR2_X1
XNOR27 STAGE26 GND STAGE27 VDD VDD GND GND NOR2_X1
XNOR28 STAGE27 GND STAGE28 VDD VDD GND GND NOR2_X1
XNOR29 STAGE28 GND STAGE29 VDD VDD GND GND NOR2_X1
XNOR30 STAGE29 GND STAGE30 VDD VDD GND GND NOR2_X1
XNOR31 STAGE30 GND STAGE31 VDD VDD GND GND NOR2_X1
XNOR32 STAGE31 GND STAGE32 VDD VDD GND GND NOR2_X1
XNOR33 STAGE32 GND STAGE33 VDD VDD GND GND NOR2_X1
XNOR34 STAGE33 GND STAGE34 VDD VDD GND GND NOR2_X1
XNOR35 STAGE34 GND STAGE35 VDD VDD GND GND NOR2_X1
XNOR36 STAGE35 GND STAGE36 VDD VDD GND GND NOR2_X1
XNOR37 STAGE36 GND STAGE37 VDD VDD GND GND NOR2_X1
XNOR38 STAGE37 GND STAGE38 VDD VDD GND GND NOR2_X1
XNOR39 STAGE38 GND STAGE39 VDD VDD GND GND NOR2_X1
XNOR40 STAGE39 GND STAGE40 VDD VDD GND GND NOR2_X1
XNOR41 STAGE40 GND STAGE41 VDD VDD GND GND NOR2_X1
XNOR42 STAGE41 GND STAGE42 VDD VDD GND GND NOR2_X1
XNOR43 STAGE42 GND STAGE43 VDD VDD GND GND NOR2_X1
XNOR44 STAGE43 GND STAGE44 VDD VDD GND GND NOR2_X1
XNOR45 STAGE44 GND STAGE45 VDD VDD GND GND NOR2_X1
XNOR46 STAGE45 GND STAGE46 VDD VDD GND GND NOR2_X1
XNOR47 STAGE46 GND STAGE47 VDD VDD GND GND NOR2_X1
XNOR48 STAGE47 GND STAGE48 VDD VDD GND GND NOR2_X1
XNOR49 STAGE48 GND STAGE49 VDD VDD GND GND NOR2_X1
XNOR50 STAGE49 GND STAGE50 VDD VDD GND GND NOR2_X1
XNOR51 STAGE50 GND STAGE51 VDD VDD GND GND NOR2_X1
XNOR52 STAGE51 GND STAGE52 VDD VDD GND GND NOR2_X1
XNOR53 STAGE52 GND STAGE53 VDD VDD GND GND NOR2_X1
XNOR54 STAGE53 GND STAGE54 VDD VDD GND GND NOR2_X1
XNOR55 STAGE54 GND STAGE55 VDD VDD GND GND NOR2_X1
XNOR56 STAGE55 GND STAGE56 VDD VDD GND GND NOR2_X1
XNOR57 STAGE56 GND STAGE57 VDD VDD GND GND NOR2_X1
XNOR58 STAGE57 GND STAGE58 VDD VDD GND GND NOR2_X1
XNOR59 STAGE58 GND STAGE59 VDD VDD GND GND NOR2_X1
XNOR60 STAGE59 GND STAGE60 VDD VDD GND GND NOR2_X1
XNOR61 STAGE60 GND STAGE61 VDD VDD GND GND NOR2_X1
XNOR62 STAGE61 GND STAGE62 VDD VDD GND GND NOR2_X1
XNOR63 STAGE62 GND STAGE63 VDD VDD GND GND NOR2_X1
XNOR64 STAGE63 GND STAGE64 VDD VDD GND GND NOR2_X1
XNOR65 STAGE64 GND STAGE65 VDD VDD GND GND NOR2_X1
XNOR66 STAGE65 GND STAGE66 VDD VDD GND GND NOR2_X1
XNOR67 STAGE66 GND STAGE67 VDD VDD GND GND NOR2_X1
XNOR68 STAGE67 GND STAGE68 VDD VDD GND GND NOR2_X1
XNOR69 STAGE68 GND STAGE69 VDD VDD GND GND NOR2_X1
XNOR70 STAGE69 GND STAGE70 VDD VDD GND GND NOR2_X1
XNOR71 STAGE70 GND STAGE71 VDD VDD GND GND NOR2_X1
XNOR72 STAGE71 GND STAGE72 VDD VDD GND GND NOR2_X1
XNOR73 STAGE72 GND STAGE73 VDD VDD GND GND NOR2_X1
XNOR74 STAGE73 GND STAGE74 VDD VDD GND GND NOR2_X1
XNOR75 STAGE74 GND STAGE75 VDD VDD GND GND NOR2_X1
XNOR76 STAGE75 GND STAGE76 VDD VDD GND GND NOR2_X1
XNOR77 STAGE76 GND STAGE77 VDD VDD GND GND NOR2_X1
XNOR78 STAGE77 GND STAGE78 VDD VDD GND GND NOR2_X1
XNOR79 STAGE78 GND STAGE79 VDD VDD GND GND NOR2_X1
XNOR80 STAGE79 GND STAGE80 VDD VDD GND GND NOR2_X1
XNOR81 STAGE80 GND STAGE81 VDD VDD GND GND NOR2_X1
XNOR82 STAGE81 GND STAGE82 VDD VDD GND GND NOR2_X1
XNOR83 STAGE82 GND STAGE83 VDD VDD GND GND NOR2_X1
XNOR84 STAGE83 GND STAGE84 VDD VDD GND GND NOR2_X1
XNOR85 STAGE84 GND STAGE85 VDD VDD GND GND NOR2_X1
XNOR86 STAGE85 GND STAGE86 VDD VDD GND GND NOR2_X1
XNOR87 STAGE86 GND STAGE87 VDD VDD GND GND NOR2_X1
XNOR88 STAGE87 GND STAGE88 VDD VDD GND GND NOR2_X1
XNOR89 STAGE88 GND STAGE89 VDD VDD GND GND NOR2_X1
XNOR90 STAGE89 GND STAGE90 VDD VDD GND GND NOR2_X1
XNOR91 STAGE90 GND STAGE91 VDD VDD GND GND NOR2_X1
XNOR92 STAGE91 GND STAGE92 VDD VDD GND GND NOR2_X1
XNOR93 STAGE92 GND STAGE93 VDD VDD GND GND NOR2_X1
XNOR94 STAGE93 GND STAGE94 VDD VDD GND GND NOR2_X1
XNOR95 STAGE94 GND STAGE95 VDD VDD GND GND NOR2_X1
XNOR96 STAGE95 GND STAGE96 VDD VDD GND GND NOR2_X1
XNOR97 STAGE96 GND STAGE97 VDD VDD GND GND NOR2_X1
XNOR98 STAGE97 GND STAGE98 VDD VDD GND GND NOR2_X1
XNOR99 STAGE98 GND STAGE99 VDD VDD GND GND NOR2_X1
XNOR100 STAGE99 GND STAGE100 VDD VDD GND GND NOR2_X1
XNOR101 STAGE100 GND STAGE101 VDD VDD GND GND NOR2_X1
XNOR102 STAGE101 GND STAGE102 VDD VDD GND GND NOR2_X1
XNOR103 STAGE102 GND STAGE103 VDD VDD GND GND NOR2_X1
XNOR104 STAGE103 GND STAGE104 VDD VDD GND GND NOR2_X1
XNOR105 STAGE104 GND STAGE105 VDD VDD GND GND NOR2_X1
XNOR106 STAGE105 GND STAGE106 VDD VDD GND GND NOR2_X1
XNOR107 STAGE106 GND STAGE107 VDD VDD GND GND NOR2_X1
XNOR108 STAGE107 GND STAGE108 VDD VDD GND GND NOR2_X1
XNOR109 STAGE108 GND STAGE109 VDD VDD GND GND NOR2_X1
XNOR110 STAGE109 GND STAGE110 VDD VDD GND GND NOR2_X1
XNOR111 STAGE110 GND STAGE111 VDD VDD GND GND NOR2_X1
XNOR112 STAGE111 GND STAGE112 VDD VDD GND GND NOR2_X1
XNOR113 STAGE112 GND STAGE113 VDD VDD GND GND NOR2_X1
XNOR114 STAGE113 GND STAGE114 VDD VDD GND GND NOR2_X1
XNOR115 STAGE114 GND STAGE115 VDD VDD GND GND NOR2_X1
XNOR116 STAGE115 GND STAGE116 VDD VDD GND GND NOR2_X1
XNOR117 STAGE116 GND STAGE117 VDD VDD GND GND NOR2_X1
XNOR118 STAGE117 GND STAGE118 VDD VDD GND GND NOR2_X1
XNOR119 STAGE118 GND myout VDD VDD GND GND NOR2_X1
C_TERM myout GND 0.0779pF

.PROBE TRAN V(myin) V(STAGE1) V(STAGE2) V(STAGE3) V(STAGE4) V(STAGE5) V(STAGE6) V(STAGE7) V(STAGE8) V(STAGE9) V(STAGE10) V(STAGE11) V(STAGE12) V(STAGE13) V(STAGE14) V(STAGE15) V(STAGE16) V(STAGE17) V(STAGE18) V(STAGE19) V(STAGE20) V(STAGE21) V(STAGE22) V(STAGE23) V(STAGE24) V(STAGE25) V(STAGE26) V(STAGE27) V(STAGE28) V(STAGE29) V(STAGE30) V(STAGE31) V(STAGE32) V(STAGE33) V(STAGE34) V(STAGE35) V(STAGE36) V(STAGE37) V(STAGE38) V(STAGE39) V(STAGE40) V(STAGE41) V(STAGE42) V(STAGE43) V(STAGE44) V(STAGE45) V(STAGE46) V(STAGE47) V(STAGE48) V(STAGE49) V(STAGE50) V(STAGE51) V(STAGE52) V(STAGE53) V(STAGE54) V(STAGE55) V(STAGE56) V(STAGE57) V(STAGE58) V(STAGE59) V(STAGE60) V(STAGE61) V(STAGE62) V(STAGE63) V(STAGE64) V(STAGE65) V(STAGE66) V(STAGE67) V(STAGE68) V(STAGE69) V(STAGE70) V(STAGE71) V(STAGE72) V(STAGE73) V(STAGE74) V(STAGE75) V(STAGE76) V(STAGE77) V(STAGE78) V(STAGE79) V(STAGE80) V(STAGE81) V(STAGE82) V(STAGE83) V(STAGE84) V(STAGE85) V(STAGE86) V(STAGE87) V(STAGE88) V(STAGE89) V(STAGE90) V(STAGE91) V(STAGE92) V(STAGE93) V(STAGE94) V(STAGE95) V(STAGE96) V(STAGE97) V(STAGE98) V(STAGE99) V(STAGE100) V(STAGE101) V(STAGE102) V(STAGE103) V(STAGE104) V(STAGE105) V(STAGE106) V(STAGE107) V(STAGE108) V(STAGE109) V(STAGE110) V(STAGE111) V(STAGE112) V(STAGE113) V(STAGE114) V(STAGE115)
.TRAN 0.1ps tend
.END

* circuit: inv tree
simulator lang=spice

.PARAM pw=<sed>pw<sed>as


.LIB <path>/back_end/spice/fet.inc CMG 

* main circuit
.INCLUDE <path>/back_end/spice/cell/OR2_X1.sp
.INCLUDE <path>/back_end/spice/cell/BUF_X4.sp
.INCLUDE <path>/back_end/spice/cell/BUF_X1.sp
.INCLUDE <path>/back_end/spice/cell/CLKBUF_X2.sp

**** SPECTRE Back Annotation
.option spef='../place_and_route/or_loop_altered.spef'
****

.TEMP 25 
.OPTION
+ INGOLD=2
+ PARHIER=LOCAL
*+ POST=CSDF
+ PROBE
+ BRIEF
+ ACCURATE
+ ABSVAR=0.05
*+ DELMAX=100fs
+ dc_pivot_check=yes

* vdd
VDD VDD GND 0.8v

* circuit under test
XBUF_I1 myin BI1 VDD VDD GND GND BUF_X4
XBUF_I2 BI1 BI2 VDD VDD GND GND BUF_X4
XBUF_I3 BI2 BI3 VDD VDD GND GND BUF_X4

XOR BI3 n_5 OR1 VDD VDD GND GND OR2_X1

XBUF_FB1 OR1 FB1 VDD VDD GND GND BUF_X4
XBUF_FB2 FB1 FB2 VDD VDD GND GND BUF_X4
XBUF_FB3 FB2 FB3 VDD VDD GND GND BUF_X4
XBUF_FB4 FB3 FB4 VDD VDD GND GND BUF_X4
XBUF_FB5 FB4 FB5 VDD VDD GND GND BUF_X4
XBUF_FB6 FB5 FB6 VDD VDD GND GND BUF_X4
XBUF_FB7 FB6 FB7 VDD VDD GND GND BUF_X4
XBUF_FB8 FB7 FB8 VDD VDD GND GND BUF_X4
XBUF_FB9 FB8 FB9 VDD VDD GND GND BUF_X4

XBUF_FB10 FB9 FB10 VDD VDD GND GND BUF_X4
XBUF_FB11 FB10 FB11 VDD VDD GND GND BUF_X4
XBUF_FB12 FB11 FB12 VDD VDD GND GND BUF_X4
XBUF_FB13 FB12 FB13 VDD VDD GND GND BUF_X4
XBUF_FB14 FB13 FB14 VDD VDD GND GND BUF_X4
XBUF_FB15 FB14 FB15 VDD VDD GND GND BUF_X4
XBUF_FB16 FB15 FB16 VDD VDD GND GND BUF_X4
XBUF_FB17 FB16 FB17 VDD VDD GND GND BUF_X4
XBUF_FB18 FB17 FB18 VDD VDD GND GND BUF_X4
XBUF_FB19 FB18 FB19 VDD VDD GND GND BUF_X4

XBUF_FB20 FB19 FB20 VDD VDD GND GND BUF_X4
XBUF_FB21 FB20 FB21 VDD VDD GND GND BUF_X4
XBUF_FB22 FB21 FB22 VDD VDD GND GND BUF_X4
XBUF_FB23 FB22 FB23 VDD VDD GND GND BUF_X4
XBUF_FB24 FB23 FB24 VDD VDD GND GND BUF_X4
XBUF_FB25 FB24 FB25 VDD VDD GND GND BUF_X4
XBUF_FB26 FB25 FB26 VDD VDD GND GND BUF_X4
XBUF_FB27 FB26 FB27 VDD VDD GND GND BUF_X4
XBUF_FB28 FB27 FB28 VDD VDD GND GND BUF_X4
XBUF_FB29 FB28 FB29 VDD VDD GND GND BUF_X4

Xcdn_loop_breaker FB29 n_5 VDD VDD GND GND CLKBUF_X2

XBUF_HT OR1 HT1 VDD VDD GND GND BUF_X1
XBUF_O1 HT1 BO1 VDD VDD GND GND BUF_X4
XBUF_O2 BO1 BO2 VDD VDD GND GND BUF_X4
XBUF_O3 BO2 myout VDD VDD GND GND BUF_X4

VIN myin 0 PULSE(0 0.8 50ps 1fs 1fs pw 20ns)

.PROBE TRAN v(myin) v(BI*) v(OR1) v(FB*) v(HT1) v(BO*) v(myout)
.NODESET OR1=0 
.TRAN 0.01PS 4000ps

.END

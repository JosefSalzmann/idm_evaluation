* circuit: cgate_test
simulator lang=spice

*.PARAM pw=<sed>pw<sed>as
.PARAM supp=0.8V slope=0.1fs
.PARAM t_init0=0.1ns t_init1=0.174ns
.PARAM baseVal=0V peakVal=0.8V tend=8100.0ns


.LIB /home/s11777724/involution_tool_library_files/backend/spice/fet.inc CMG

* main circuit
.INCLUDE /home/s11777724/involution_tool_library_files/backend/spice/cell/BUF_X8.sp
.INCLUDE cgate.sp

**** SPECTRE Back Annotation
.option spef='/home/s11777724/JS/idm_evaluation/cgate_test/place_and_route/cgate_test_restitch.spef'
****

.TEMP 25
.OPTION
+ INGOLD=2
+ PARHIER=LOCAL
*+ POST=CSDF
+ PROBE
+ BRIEF
+ ACCURATE
+ ABSVAR=0.0001
+ DVDT=2
+ RELTOL=1e-11
*+ DELMAX=100fs
+ dc_pivot_check=yes

* vdd
VDD VDD GND 0.8v

.PARAM t_a_0=10ns
.PARAM t_a_1=13.333333ns
.PARAM t_a_2=15ns
.PARAM t_a_3=18.333333ns
.PARAM t_a_4=20ns
.PARAM t_a_5=23.333333ns
.PARAM t_a_6=25ns
.PARAM t_a_7=28.333333ns
.PARAM t_a_8=30ns
.PARAM t_a_9=33.333333ns
.PARAM t_a_10=35ns
.PARAM t_a_11=38.333333ns
.PARAM t_a_12=40ns
.PARAM t_a_13=43.333333ns
.PARAM t_a_14=45ns
.PARAM t_a_15=48.333333ns
.PARAM t_a_16=50ns
.PARAM t_a_17=53.333333ns
.PARAM t_a_18=55ns
.PARAM t_a_19=58.333333ns
.PARAM t_a_20=60ns
.PARAM t_a_21=63.333333ns
.PARAM t_a_22=65ns
.PARAM t_a_23=68.333333ns
.PARAM t_a_24=70ns
.PARAM t_a_25=73.333333ns
.PARAM t_a_26=75ns
.PARAM t_a_27=78.333333ns
.PARAM t_a_28=80ns
.PARAM t_a_29=83.333333ns
.PARAM t_a_30=85ns
.PARAM t_a_31=88.333333ns
.PARAM t_a_32=90ns
.PARAM t_a_33=93.333333ns
.PARAM t_a_34=95ns
.PARAM t_a_35=98.333333ns
.PARAM t_a_36=100ns
.PARAM t_a_37=103.333333ns
.PARAM t_a_38=105ns
.PARAM t_a_39=108.333333ns
.PARAM t_a_40=110ns
.PARAM t_a_41=113.333333ns
.PARAM t_a_42=115ns
.PARAM t_a_43=118.333333ns
.PARAM t_a_44=120ns
.PARAM t_a_45=123.333333ns
.PARAM t_a_46=125ns
.PARAM t_a_47=128.333333ns
.PARAM t_a_48=130ns
.PARAM t_a_49=133.333333ns
.PARAM t_a_50=135ns
.PARAM t_a_51=138.333333ns
.PARAM t_a_52=140ns
.PARAM t_a_53=143.333333ns
.PARAM t_a_54=145ns
.PARAM t_a_55=148.333333ns
.PARAM t_a_56=150ns
.PARAM t_a_57=153.333333ns
.PARAM t_a_58=155ns
.PARAM t_a_59=158.333333ns
.PARAM t_a_60=160ns
.PARAM t_a_61=163.333333ns
.PARAM t_a_62=165ns
.PARAM t_a_63=168.333333ns
.PARAM t_a_64=170ns
.PARAM t_a_65=173.333333ns
.PARAM t_a_66=175ns
.PARAM t_a_67=178.333333ns
.PARAM t_a_68=180ns
.PARAM t_a_69=183.333333ns
.PARAM t_a_70=185ns
.PARAM t_a_71=188.333333ns
.PARAM t_a_72=190ns
.PARAM t_a_73=193.333333ns
.PARAM t_a_74=195ns
.PARAM t_a_75=198.333333ns
.PARAM t_a_76=200ns
.PARAM t_a_77=203.333333ns
.PARAM t_a_78=205ns
.PARAM t_a_79=208.333333ns
.PARAM t_a_80=210ns
.PARAM t_a_81=213.333333ns
.PARAM t_a_82=215ns
.PARAM t_a_83=218.333333ns
.PARAM t_a_84=220ns
.PARAM t_a_85=223.333333ns
.PARAM t_a_86=225ns
.PARAM t_a_87=228.333333ns
.PARAM t_a_88=230ns
.PARAM t_a_89=233.333333ns
.PARAM t_a_90=235ns
.PARAM t_a_91=238.333333ns
.PARAM t_a_92=240ns
.PARAM t_a_93=243.333333ns
.PARAM t_a_94=245ns
.PARAM t_a_95=248.333333ns
.PARAM t_a_96=250ns
.PARAM t_a_97=253.333333ns
.PARAM t_a_98=255ns
.PARAM t_a_99=258.333333ns
.PARAM t_a_100=260ns
.PARAM t_a_101=263.333333ns
.PARAM t_a_102=265ns
.PARAM t_a_103=268.333333ns
.PARAM t_a_104=270ns
.PARAM t_a_105=273.333333ns
.PARAM t_a_106=275ns
.PARAM t_a_107=278.333333ns
.PARAM t_a_108=280ns
.PARAM t_a_109=283.333333ns
.PARAM t_a_110=285ns
.PARAM t_a_111=288.333333ns
.PARAM t_a_112=290ns
.PARAM t_a_113=293.333333ns
.PARAM t_a_114=295ns
.PARAM t_a_115=298.333333ns
.PARAM t_a_116=300ns
.PARAM t_a_117=303.333333ns
.PARAM t_a_118=305ns
.PARAM t_a_119=308.333333ns
.PARAM t_a_120=310ns
.PARAM t_a_121=313.333333ns
.PARAM t_a_122=315ns
.PARAM t_a_123=318.333333ns
.PARAM t_a_124=320ns
.PARAM t_a_125=323.333333ns
.PARAM t_a_126=325ns
.PARAM t_a_127=328.333333ns
.PARAM t_a_128=330ns
.PARAM t_a_129=333.333333ns
.PARAM t_a_130=335ns
.PARAM t_a_131=338.333333ns
.PARAM t_a_132=340ns
.PARAM t_a_133=343.333333ns
.PARAM t_a_134=345ns
.PARAM t_a_135=348.333333ns
.PARAM t_a_136=350ns
.PARAM t_a_137=353.333333ns
.PARAM t_a_138=355ns
.PARAM t_a_139=358.333333ns
.PARAM t_a_140=360ns
.PARAM t_a_141=363.333333ns
.PARAM t_a_142=365ns
.PARAM t_a_143=368.333333ns
.PARAM t_a_144=370ns
.PARAM t_a_145=373.333333ns
.PARAM t_a_146=375ns
.PARAM t_a_147=378.333333ns
.PARAM t_a_148=380ns
.PARAM t_a_149=383.333333ns
.PARAM t_a_150=385ns
.PARAM t_a_151=388.333333ns
.PARAM t_a_152=390ns
.PARAM t_a_153=393.333333ns
.PARAM t_a_154=395ns
.PARAM t_a_155=398.333333ns
.PARAM t_a_156=400ns
.PARAM t_a_157=403.333333ns
.PARAM t_a_158=405ns
.PARAM t_a_159=408.333333ns
.PARAM t_a_160=410ns
.PARAM t_a_161=413.333333ns
.PARAM t_a_162=415ns
.PARAM t_a_163=418.333333ns
.PARAM t_a_164=420ns
.PARAM t_a_165=423.333333ns
.PARAM t_a_166=425ns
.PARAM t_a_167=428.333333ns
.PARAM t_a_168=430ns
.PARAM t_a_169=433.333333ns
.PARAM t_a_170=435ns
.PARAM t_a_171=438.333333ns
.PARAM t_a_172=440ns
.PARAM t_a_173=443.333333ns
.PARAM t_a_174=445ns
.PARAM t_a_175=448.333333ns
.PARAM t_a_176=450ns
.PARAM t_a_177=453.333333ns
.PARAM t_a_178=455ns
.PARAM t_a_179=458.333333ns
.PARAM t_a_180=460ns
.PARAM t_a_181=463.333333ns
.PARAM t_a_182=465ns
.PARAM t_a_183=468.333333ns
.PARAM t_a_184=470ns
.PARAM t_a_185=473.333333ns
.PARAM t_a_186=475ns
.PARAM t_a_187=478.333333ns
.PARAM t_a_188=480ns
.PARAM t_a_189=483.333333ns
.PARAM t_a_190=485ns
.PARAM t_a_191=488.333333ns
.PARAM t_a_192=490ns
.PARAM t_a_193=493.333333ns
.PARAM t_a_194=495ns
.PARAM t_a_195=498.333333ns
.PARAM t_a_196=500ns
.PARAM t_a_197=503.333333ns
.PARAM t_a_198=505ns
.PARAM t_a_199=508.333333ns
.PARAM t_a_200=510ns
.PARAM t_a_201=513.333333ns
.PARAM t_a_202=515ns
.PARAM t_a_203=518.333333ns
.PARAM t_a_204=520ns
.PARAM t_a_205=523.333333ns
.PARAM t_a_206=525ns
.PARAM t_a_207=528.333333ns
.PARAM t_a_208=530ns
.PARAM t_a_209=533.333333ns
.PARAM t_a_210=535ns
.PARAM t_a_211=538.333333ns
.PARAM t_a_212=540ns
.PARAM t_a_213=543.333333ns
.PARAM t_a_214=545ns
.PARAM t_a_215=548.333333ns
.PARAM t_a_216=550ns
.PARAM t_a_217=553.333333ns
.PARAM t_a_218=555ns
.PARAM t_a_219=558.333333ns
.PARAM t_a_220=560ns
.PARAM t_a_221=563.333333ns
.PARAM t_a_222=565ns
.PARAM t_a_223=568.333333ns
.PARAM t_a_224=570ns
.PARAM t_a_225=573.333333ns
.PARAM t_a_226=575ns
.PARAM t_a_227=578.333333ns
.PARAM t_a_228=580ns
.PARAM t_a_229=583.333333ns
.PARAM t_a_230=585ns
.PARAM t_a_231=588.333333ns
.PARAM t_a_232=590ns
.PARAM t_a_233=593.333333ns
.PARAM t_a_234=595ns
.PARAM t_a_235=598.333333ns
.PARAM t_a_236=600ns
.PARAM t_a_237=603.333333ns
.PARAM t_a_238=605ns
.PARAM t_a_239=608.333333ns
.PARAM t_a_240=610ns
.PARAM t_a_241=613.333333ns
.PARAM t_a_242=615ns
.PARAM t_a_243=618.333333ns
.PARAM t_a_244=620ns
.PARAM t_a_245=623.333333ns
.PARAM t_a_246=625ns
.PARAM t_a_247=628.333333ns
.PARAM t_a_248=630ns
.PARAM t_a_249=633.333333ns
.PARAM t_a_250=635ns
.PARAM t_a_251=638.333333ns
.PARAM t_a_252=640ns
.PARAM t_a_253=643.333333ns
.PARAM t_a_254=645ns
.PARAM t_a_255=648.333333ns
.PARAM t_a_256=650ns
.PARAM t_a_257=653.333333ns
.PARAM t_a_258=655ns
.PARAM t_a_259=658.333333ns
.PARAM t_a_260=660ns
.PARAM t_a_261=663.333333ns
.PARAM t_a_262=665ns
.PARAM t_a_263=668.333333ns
.PARAM t_a_264=670ns
.PARAM t_a_265=673.333333ns
.PARAM t_a_266=675ns
.PARAM t_a_267=678.333333ns
.PARAM t_a_268=680ns
.PARAM t_a_269=683.333333ns
.PARAM t_a_270=685ns
.PARAM t_a_271=688.333333ns
.PARAM t_a_272=690ns
.PARAM t_a_273=693.333333ns
.PARAM t_a_274=695ns
.PARAM t_a_275=698.333333ns
.PARAM t_a_276=700ns
.PARAM t_a_277=703.333333ns
.PARAM t_a_278=705ns
.PARAM t_a_279=708.333333ns
.PARAM t_a_280=710ns
.PARAM t_a_281=713.333333ns
.PARAM t_a_282=715ns
.PARAM t_a_283=718.333333ns
.PARAM t_a_284=720ns
.PARAM t_a_285=723.333333ns
.PARAM t_a_286=725ns
.PARAM t_a_287=728.333333ns
.PARAM t_a_288=730ns
.PARAM t_a_289=733.333333ns
.PARAM t_a_290=735ns
.PARAM t_a_291=738.333333ns
.PARAM t_a_292=740ns
.PARAM t_a_293=743.333333ns
.PARAM t_a_294=745ns
.PARAM t_a_295=748.333333ns
.PARAM t_a_296=750ns
.PARAM t_a_297=753.333333ns
.PARAM t_a_298=755ns
.PARAM t_a_299=758.333333ns
.PARAM t_a_300=760ns
.PARAM t_a_301=763.333333ns
.PARAM t_a_302=765ns
.PARAM t_a_303=768.333333ns
.PARAM t_a_304=770ns
.PARAM t_a_305=773.333333ns
.PARAM t_a_306=775ns
.PARAM t_a_307=778.333333ns
.PARAM t_a_308=780ns
.PARAM t_a_309=783.333333ns
.PARAM t_a_310=785ns
.PARAM t_a_311=788.333333ns
.PARAM t_a_312=790ns
.PARAM t_a_313=793.333333ns
.PARAM t_a_314=795ns
.PARAM t_a_315=798.333333ns
.PARAM t_a_316=800ns
.PARAM t_a_317=803.333333ns
.PARAM t_a_318=805ns
.PARAM t_a_319=808.333333ns
.PARAM t_a_320=810ns
.PARAM t_a_321=813.333333ns
.PARAM t_a_322=815ns
.PARAM t_a_323=818.333333ns
.PARAM t_a_324=820ns
.PARAM t_a_325=823.333333ns
.PARAM t_a_326=825ns
.PARAM t_a_327=828.333333ns
.PARAM t_a_328=830ns
.PARAM t_a_329=833.333333ns
.PARAM t_a_330=835ns
.PARAM t_a_331=838.333333ns
.PARAM t_a_332=840ns
.PARAM t_a_333=843.333333ns
.PARAM t_a_334=845ns
.PARAM t_a_335=848.333333ns
.PARAM t_a_336=850ns
.PARAM t_a_337=853.333333ns
.PARAM t_a_338=855ns
.PARAM t_a_339=858.333333ns
.PARAM t_a_340=860ns
.PARAM t_a_341=863.333333ns
.PARAM t_a_342=865ns
.PARAM t_a_343=868.333333ns
.PARAM t_a_344=870ns
.PARAM t_a_345=873.333333ns
.PARAM t_a_346=875ns
.PARAM t_a_347=878.333333ns
.PARAM t_a_348=880ns
.PARAM t_a_349=883.333333ns
.PARAM t_a_350=885ns
.PARAM t_a_351=888.333333ns
.PARAM t_a_352=890ns
.PARAM t_a_353=893.333333ns
.PARAM t_a_354=895ns
.PARAM t_a_355=898.333333ns
.PARAM t_a_356=900ns
.PARAM t_a_357=903.333333ns
.PARAM t_a_358=905ns
.PARAM t_a_359=908.333333ns
.PARAM t_a_360=910ns
.PARAM t_a_361=913.333333ns
.PARAM t_a_362=915ns
.PARAM t_a_363=918.333333ns
.PARAM t_a_364=920ns
.PARAM t_a_365=923.333333ns
.PARAM t_a_366=925ns
.PARAM t_a_367=928.333333ns
.PARAM t_a_368=930ns
.PARAM t_a_369=933.333333ns
.PARAM t_a_370=935ns
.PARAM t_a_371=938.333333ns
.PARAM t_a_372=940ns
.PARAM t_a_373=943.333333ns
.PARAM t_a_374=945ns
.PARAM t_a_375=948.333333ns
.PARAM t_a_376=950ns
.PARAM t_a_377=953.333333ns
.PARAM t_a_378=955ns
.PARAM t_a_379=958.333333ns
.PARAM t_a_380=960ns
.PARAM t_a_381=963.333333ns
.PARAM t_a_382=965ns
.PARAM t_a_383=968.333333ns
.PARAM t_a_384=970ns
.PARAM t_a_385=973.333333ns
.PARAM t_a_386=975ns
.PARAM t_a_387=978.333333ns
.PARAM t_a_388=980ns
.PARAM t_a_389=983.333333ns
.PARAM t_a_390=985ns
.PARAM t_a_391=988.333333ns
.PARAM t_a_392=990ns
.PARAM t_a_393=993.333333ns
.PARAM t_a_394=995ns
.PARAM t_a_395=998.333333ns
.PARAM t_a_396=1000ns
.PARAM t_a_397=1003.333333ns
.PARAM t_a_398=1005ns
.PARAM t_a_399=1008.333333ns
.PARAM t_a_400=1010ns
.PARAM t_a_401=1013.333333ns
.PARAM t_a_402=1015ns
.PARAM t_a_403=1018.333333ns
.PARAM t_a_404=1020ns
.PARAM t_a_405=1023.333333ns
.PARAM t_a_406=1025ns
.PARAM t_a_407=1028.333333ns
.PARAM t_a_408=1030ns
.PARAM t_a_409=1033.333333ns
.PARAM t_a_410=1035ns
.PARAM t_a_411=1038.333333ns
.PARAM t_a_412=1040ns
.PARAM t_a_413=1043.333333ns
.PARAM t_a_414=1045ns
.PARAM t_a_415=1048.333333ns
.PARAM t_a_416=1050ns
.PARAM t_a_417=1053.333333ns
.PARAM t_a_418=1055ns
.PARAM t_a_419=1058.333333ns
.PARAM t_a_420=1060ns
.PARAM t_a_421=1063.333333ns
.PARAM t_a_422=1065ns
.PARAM t_a_423=1068.333333ns
.PARAM t_a_424=1070ns
.PARAM t_a_425=1073.333333ns
.PARAM t_a_426=1075ns
.PARAM t_a_427=1078.333333ns
.PARAM t_a_428=1080ns
.PARAM t_a_429=1083.333333ns
.PARAM t_a_430=1085ns
.PARAM t_a_431=1088.333333ns
.PARAM t_a_432=1090ns
.PARAM t_a_433=1093.333333ns
.PARAM t_a_434=1095ns
.PARAM t_a_435=1098.333333ns
.PARAM t_a_436=1100ns
.PARAM t_a_437=1103.333333ns
.PARAM t_a_438=1105ns
.PARAM t_a_439=1108.333333ns
.PARAM t_a_440=1110ns
.PARAM t_a_441=1113.333333ns
.PARAM t_a_442=1115ns
.PARAM t_a_443=1118.333333ns
.PARAM t_a_444=1120ns
.PARAM t_a_445=1123.333333ns
.PARAM t_a_446=1125ns
.PARAM t_a_447=1128.333333ns
.PARAM t_a_448=1130ns
.PARAM t_a_449=1133.333333ns
.PARAM t_a_450=1135ns
.PARAM t_a_451=1138.333333ns
.PARAM t_a_452=1140ns
.PARAM t_a_453=1143.333333ns
.PARAM t_a_454=1145ns
.PARAM t_a_455=1148.333333ns
.PARAM t_a_456=1150ns
.PARAM t_a_457=1153.333333ns
.PARAM t_a_458=1155ns
.PARAM t_a_459=1158.333333ns
.PARAM t_a_460=1160ns
.PARAM t_a_461=1163.333333ns
.PARAM t_a_462=1165ns
.PARAM t_a_463=1168.333333ns
.PARAM t_a_464=1170ns
.PARAM t_a_465=1173.333333ns
.PARAM t_a_466=1175ns
.PARAM t_a_467=1178.333333ns
.PARAM t_a_468=1180ns
.PARAM t_a_469=1183.333333ns
.PARAM t_a_470=1185ns
.PARAM t_a_471=1188.333333ns
.PARAM t_a_472=1190ns
.PARAM t_a_473=1193.333333ns
.PARAM t_a_474=1195ns
.PARAM t_a_475=1198.333333ns
.PARAM t_a_476=1200ns
.PARAM t_a_477=1203.333333ns
.PARAM t_a_478=1205ns
.PARAM t_a_479=1208.333333ns
.PARAM t_a_480=1210ns
.PARAM t_a_481=1213.333333ns
.PARAM t_a_482=1215ns
.PARAM t_a_483=1218.333333ns
.PARAM t_a_484=1220ns
.PARAM t_a_485=1223.333333ns
.PARAM t_a_486=1225ns
.PARAM t_a_487=1228.333333ns
.PARAM t_a_488=1230ns
.PARAM t_a_489=1233.333333ns
.PARAM t_a_490=1235ns
.PARAM t_a_491=1238.333333ns
.PARAM t_a_492=1240ns
.PARAM t_a_493=1243.333333ns
.PARAM t_a_494=1245ns
.PARAM t_a_495=1248.333333ns
.PARAM t_a_496=1250ns
.PARAM t_a_497=1253.333333ns
.PARAM t_a_498=1255ns
.PARAM t_a_499=1258.333333ns
.PARAM t_a_500=1260ns
.PARAM t_a_501=1263.333333ns
.PARAM t_a_502=1265ns
.PARAM t_a_503=1268.333333ns
.PARAM t_a_504=1270ns
.PARAM t_a_505=1273.333333ns
.PARAM t_a_506=1275ns
.PARAM t_a_507=1278.333333ns
.PARAM t_a_508=1280ns
.PARAM t_a_509=1283.333333ns
.PARAM t_a_510=1285ns
.PARAM t_a_511=1288.333333ns
.PARAM t_a_512=1290ns
.PARAM t_a_513=1293.333333ns
.PARAM t_a_514=1295ns
.PARAM t_a_515=1298.333333ns
.PARAM t_a_516=1300ns
.PARAM t_a_517=1303.333333ns
.PARAM t_a_518=1305ns
.PARAM t_a_519=1308.333333ns
.PARAM t_a_520=1310ns
.PARAM t_a_521=1313.333333ns
.PARAM t_a_522=1315ns
.PARAM t_a_523=1318.333333ns
.PARAM t_a_524=1320ns
.PARAM t_a_525=1323.333333ns
.PARAM t_a_526=1325ns
.PARAM t_a_527=1328.333333ns
.PARAM t_a_528=1330ns
.PARAM t_a_529=1333.333333ns
.PARAM t_a_530=1335ns
.PARAM t_a_531=1338.333333ns
.PARAM t_a_532=1340ns
.PARAM t_a_533=1343.333333ns
.PARAM t_a_534=1345ns
.PARAM t_a_535=1348.333333ns
.PARAM t_a_536=1350ns
.PARAM t_a_537=1353.333333ns
.PARAM t_a_538=1355ns
.PARAM t_a_539=1358.333333ns
.PARAM t_a_540=1360ns
.PARAM t_a_541=1363.333333ns
.PARAM t_a_542=1365ns
.PARAM t_a_543=1368.333333ns
.PARAM t_a_544=1370ns
.PARAM t_a_545=1373.333333ns
.PARAM t_a_546=1375ns
.PARAM t_a_547=1378.333333ns
.PARAM t_a_548=1380ns
.PARAM t_a_549=1383.333333ns
.PARAM t_a_550=1385ns
.PARAM t_a_551=1388.333333ns
.PARAM t_a_552=1390ns
.PARAM t_a_553=1393.333333ns
.PARAM t_a_554=1395ns
.PARAM t_a_555=1398.333333ns
.PARAM t_a_556=1400ns
.PARAM t_a_557=1403.333333ns
.PARAM t_a_558=1405ns
.PARAM t_a_559=1408.333333ns
.PARAM t_a_560=1410ns
.PARAM t_a_561=1413.333333ns
.PARAM t_a_562=1415ns
.PARAM t_a_563=1418.333333ns
.PARAM t_a_564=1420ns
.PARAM t_a_565=1423.333333ns
.PARAM t_a_566=1425ns
.PARAM t_a_567=1428.333333ns
.PARAM t_a_568=1430ns
.PARAM t_a_569=1433.333333ns
.PARAM t_a_570=1435ns
.PARAM t_a_571=1438.333333ns
.PARAM t_a_572=1440ns
.PARAM t_a_573=1443.333333ns
.PARAM t_a_574=1445ns
.PARAM t_a_575=1448.333333ns
.PARAM t_a_576=1450ns
.PARAM t_a_577=1453.333333ns
.PARAM t_a_578=1455ns
.PARAM t_a_579=1458.333333ns
.PARAM t_a_580=1460ns
.PARAM t_a_581=1463.333333ns
.PARAM t_a_582=1465ns
.PARAM t_a_583=1468.333333ns
.PARAM t_a_584=1470ns
.PARAM t_a_585=1473.333333ns
.PARAM t_a_586=1475ns
.PARAM t_a_587=1478.333333ns
.PARAM t_a_588=1480ns
.PARAM t_a_589=1483.333333ns
.PARAM t_a_590=1485ns
.PARAM t_a_591=1488.333333ns
.PARAM t_a_592=1490ns
.PARAM t_a_593=1493.333333ns
.PARAM t_a_594=1495ns
.PARAM t_a_595=1498.333333ns
.PARAM t_a_596=1500ns
.PARAM t_a_597=1503.333333ns
.PARAM t_a_598=1505ns
.PARAM t_a_599=1508.333333ns
.PARAM t_a_600=1510ns
.PARAM t_a_601=1513.333333ns
.PARAM t_a_602=1515ns
.PARAM t_a_603=1518.333333ns
.PARAM t_a_604=1520ns
.PARAM t_a_605=1523.333333ns
.PARAM t_a_606=1525ns
.PARAM t_a_607=1528.333333ns
.PARAM t_a_608=1530ns
.PARAM t_a_609=1533.333333ns
.PARAM t_a_610=1535ns
.PARAM t_a_611=1538.333333ns
.PARAM t_a_612=1540ns
.PARAM t_a_613=1543.333333ns
.PARAM t_a_614=1545ns
.PARAM t_a_615=1548.333333ns
.PARAM t_a_616=1550ns
.PARAM t_a_617=1553.333333ns
.PARAM t_a_618=1555ns
.PARAM t_a_619=1558.333333ns
.PARAM t_a_620=1560ns
.PARAM t_a_621=1563.333333ns
.PARAM t_a_622=1565ns
.PARAM t_a_623=1568.333333ns
.PARAM t_a_624=1570ns
.PARAM t_a_625=1573.333333ns
.PARAM t_a_626=1575ns
.PARAM t_a_627=1578.333333ns
.PARAM t_a_628=1580ns
.PARAM t_a_629=1583.333333ns
.PARAM t_a_630=1585ns
.PARAM t_a_631=1588.333333ns
.PARAM t_a_632=1590ns
.PARAM t_a_633=1593.333333ns
.PARAM t_a_634=1595ns
.PARAM t_a_635=1598.333333ns
.PARAM t_a_636=1600ns
.PARAM t_a_637=1603.333333ns
.PARAM t_a_638=1605ns
.PARAM t_a_639=1608.333333ns
.PARAM t_a_640=1610ns
.PARAM t_a_641=1613.333333ns
.PARAM t_a_642=1615ns
.PARAM t_a_643=1618.333333ns
.PARAM t_a_644=1620ns
.PARAM t_a_645=1623.333333ns
.PARAM t_a_646=1625ns
.PARAM t_a_647=1628.333333ns
.PARAM t_a_648=1630ns
.PARAM t_a_649=1633.333333ns
.PARAM t_a_650=1635ns
.PARAM t_a_651=1638.333333ns
.PARAM t_a_652=1640ns
.PARAM t_a_653=1643.333333ns
.PARAM t_a_654=1645ns
.PARAM t_a_655=1648.333333ns
.PARAM t_a_656=1650ns
.PARAM t_a_657=1653.333333ns
.PARAM t_a_658=1655ns
.PARAM t_a_659=1658.333333ns
.PARAM t_a_660=1660ns
.PARAM t_a_661=1663.333333ns
.PARAM t_a_662=1665ns
.PARAM t_a_663=1668.333333ns
.PARAM t_a_664=1670ns
.PARAM t_a_665=1673.333333ns
.PARAM t_a_666=1675ns
.PARAM t_a_667=1678.333333ns
.PARAM t_a_668=1680ns
.PARAM t_a_669=1683.333333ns
.PARAM t_a_670=1685ns
.PARAM t_a_671=1688.333333ns
.PARAM t_a_672=1690ns
.PARAM t_a_673=1693.333333ns
.PARAM t_a_674=1695ns
.PARAM t_a_675=1698.333333ns
.PARAM t_a_676=1700ns
.PARAM t_a_677=1703.333333ns
.PARAM t_a_678=1705ns
.PARAM t_a_679=1708.333333ns
.PARAM t_a_680=1710ns
.PARAM t_a_681=1713.333333ns
.PARAM t_a_682=1715ns
.PARAM t_a_683=1718.333333ns
.PARAM t_a_684=1720ns
.PARAM t_a_685=1723.333333ns
.PARAM t_a_686=1725ns
.PARAM t_a_687=1728.333333ns
.PARAM t_a_688=1730ns
.PARAM t_a_689=1733.333333ns
.PARAM t_a_690=1735ns
.PARAM t_a_691=1738.333333ns
.PARAM t_a_692=1740ns
.PARAM t_a_693=1743.333333ns
.PARAM t_a_694=1745ns
.PARAM t_a_695=1748.333333ns
.PARAM t_a_696=1750ns
.PARAM t_a_697=1753.333333ns
.PARAM t_a_698=1755ns
.PARAM t_a_699=1758.333333ns
.PARAM t_a_700=1760ns
.PARAM t_a_701=1763.333333ns
.PARAM t_a_702=1765ns
.PARAM t_a_703=1768.333333ns
.PARAM t_a_704=1770ns
.PARAM t_a_705=1773.333333ns
.PARAM t_a_706=1775ns
.PARAM t_a_707=1778.333333ns
.PARAM t_a_708=1780ns
.PARAM t_a_709=1783.333333ns
.PARAM t_a_710=1785ns
.PARAM t_a_711=1788.333333ns
.PARAM t_a_712=1790ns
.PARAM t_a_713=1793.333333ns
.PARAM t_a_714=1795ns
.PARAM t_a_715=1798.333333ns
.PARAM t_a_716=1800ns
.PARAM t_a_717=1803.333333ns
.PARAM t_a_718=1805ns
.PARAM t_a_719=1808.333333ns
.PARAM t_a_720=1810ns
.PARAM t_a_721=1813.333333ns
.PARAM t_a_722=1815ns
.PARAM t_a_723=1818.333333ns
.PARAM t_a_724=1820ns
.PARAM t_a_725=1823.333333ns
.PARAM t_a_726=1825ns
.PARAM t_a_727=1828.333333ns
.PARAM t_a_728=1830ns
.PARAM t_a_729=1833.333333ns
.PARAM t_a_730=1835ns
.PARAM t_a_731=1838.333333ns
.PARAM t_a_732=1840ns
.PARAM t_a_733=1843.333333ns
.PARAM t_a_734=1845ns
.PARAM t_a_735=1848.333333ns
.PARAM t_a_736=1850ns
.PARAM t_a_737=1853.333333ns
.PARAM t_a_738=1855ns
.PARAM t_a_739=1858.333333ns
.PARAM t_a_740=1860ns
.PARAM t_a_741=1863.333333ns
.PARAM t_a_742=1865ns
.PARAM t_a_743=1868.333333ns
.PARAM t_a_744=1870ns
.PARAM t_a_745=1873.333333ns
.PARAM t_a_746=1875ns
.PARAM t_a_747=1878.333333ns
.PARAM t_a_748=1880ns
.PARAM t_a_749=1883.333333ns
.PARAM t_a_750=1885ns
.PARAM t_a_751=1888.333333ns
.PARAM t_a_752=1890ns
.PARAM t_a_753=1893.333333ns
.PARAM t_a_754=1895ns
.PARAM t_a_755=1898.333333ns
.PARAM t_a_756=1900ns
.PARAM t_a_757=1903.333333ns
.PARAM t_a_758=1905ns
.PARAM t_a_759=1908.333333ns
.PARAM t_a_760=1910ns
.PARAM t_a_761=1913.333333ns
.PARAM t_a_762=1915ns
.PARAM t_a_763=1918.333333ns
.PARAM t_a_764=1920ns
.PARAM t_a_765=1923.333333ns
.PARAM t_a_766=1925ns
.PARAM t_a_767=1928.333333ns
.PARAM t_a_768=1930ns
.PARAM t_a_769=1933.333333ns
.PARAM t_a_770=1935ns
.PARAM t_a_771=1938.333333ns
.PARAM t_a_772=1940ns
.PARAM t_a_773=1943.333333ns
.PARAM t_a_774=1945ns
.PARAM t_a_775=1948.333333ns
.PARAM t_a_776=1950ns
.PARAM t_a_777=1953.333333ns
.PARAM t_a_778=1955ns
.PARAM t_a_779=1958.333333ns
.PARAM t_a_780=1960ns
.PARAM t_a_781=1963.333333ns
.PARAM t_a_782=1965ns
.PARAM t_a_783=1968.333333ns
.PARAM t_a_784=1970ns
.PARAM t_a_785=1973.333333ns
.PARAM t_a_786=1975ns
.PARAM t_a_787=1978.333333ns
.PARAM t_a_788=1980ns
.PARAM t_a_789=1983.333333ns
.PARAM t_a_790=1985ns
.PARAM t_a_791=1988.333333ns
.PARAM t_a_792=1990ns
.PARAM t_a_793=1993.333333ns
.PARAM t_a_794=1995ns
.PARAM t_a_795=1998.333333ns
.PARAM t_a_796=2000ns
.PARAM t_a_797=2003.333333ns
.PARAM t_a_798=2005ns
.PARAM t_a_799=2008.333333ns
.PARAM t_b_0=9.8ns
.PARAM t_b_1=11.666667ns
.PARAM t_b_2=14.801ns
.PARAM t_b_3=16.666667ns
.PARAM t_b_4=19.802ns
.PARAM t_b_5=21.666667ns
.PARAM t_b_6=24.803ns
.PARAM t_b_7=26.666667ns
.PARAM t_b_8=29.804ns
.PARAM t_b_9=31.666667ns
.PARAM t_b_10=34.805ns
.PARAM t_b_11=36.666667ns
.PARAM t_b_12=39.806ns
.PARAM t_b_13=41.666667ns
.PARAM t_b_14=44.807ns
.PARAM t_b_15=46.666667ns
.PARAM t_b_16=49.808ns
.PARAM t_b_17=51.666667ns
.PARAM t_b_18=54.809ns
.PARAM t_b_19=56.666667ns
.PARAM t_b_20=59.81ns
.PARAM t_b_21=61.666667ns
.PARAM t_b_22=64.811ns
.PARAM t_b_23=66.666667ns
.PARAM t_b_24=69.812ns
.PARAM t_b_25=71.666667ns
.PARAM t_b_26=74.813ns
.PARAM t_b_27=76.666667ns
.PARAM t_b_28=79.814ns
.PARAM t_b_29=81.666667ns
.PARAM t_b_30=84.815ns
.PARAM t_b_31=86.666667ns
.PARAM t_b_32=89.816ns
.PARAM t_b_33=91.666667ns
.PARAM t_b_34=94.817ns
.PARAM t_b_35=96.666667ns
.PARAM t_b_36=99.818ns
.PARAM t_b_37=101.666667ns
.PARAM t_b_38=104.819ns
.PARAM t_b_39=106.666667ns
.PARAM t_b_40=109.82ns
.PARAM t_b_41=111.666667ns
.PARAM t_b_42=114.821ns
.PARAM t_b_43=116.666667ns
.PARAM t_b_44=119.822ns
.PARAM t_b_45=121.666667ns
.PARAM t_b_46=124.823ns
.PARAM t_b_47=126.666667ns
.PARAM t_b_48=129.824ns
.PARAM t_b_49=131.666667ns
.PARAM t_b_50=134.825ns
.PARAM t_b_51=136.666667ns
.PARAM t_b_52=139.826ns
.PARAM t_b_53=141.666667ns
.PARAM t_b_54=144.827ns
.PARAM t_b_55=146.666667ns
.PARAM t_b_56=149.828ns
.PARAM t_b_57=151.666667ns
.PARAM t_b_58=154.829ns
.PARAM t_b_59=156.666667ns
.PARAM t_b_60=159.83ns
.PARAM t_b_61=161.666667ns
.PARAM t_b_62=164.831ns
.PARAM t_b_63=166.666667ns
.PARAM t_b_64=169.832ns
.PARAM t_b_65=171.666667ns
.PARAM t_b_66=174.833ns
.PARAM t_b_67=176.666667ns
.PARAM t_b_68=179.834ns
.PARAM t_b_69=181.666667ns
.PARAM t_b_70=184.835ns
.PARAM t_b_71=186.666667ns
.PARAM t_b_72=189.836ns
.PARAM t_b_73=191.666667ns
.PARAM t_b_74=194.837ns
.PARAM t_b_75=196.666667ns
.PARAM t_b_76=199.838ns
.PARAM t_b_77=201.666667ns
.PARAM t_b_78=204.839ns
.PARAM t_b_79=206.666667ns
.PARAM t_b_80=209.84ns
.PARAM t_b_81=211.666667ns
.PARAM t_b_82=214.841ns
.PARAM t_b_83=216.666667ns
.PARAM t_b_84=219.842ns
.PARAM t_b_85=221.666667ns
.PARAM t_b_86=224.843ns
.PARAM t_b_87=226.666667ns
.PARAM t_b_88=229.844ns
.PARAM t_b_89=231.666667ns
.PARAM t_b_90=234.845ns
.PARAM t_b_91=236.666667ns
.PARAM t_b_92=239.846ns
.PARAM t_b_93=241.666667ns
.PARAM t_b_94=244.847ns
.PARAM t_b_95=246.666667ns
.PARAM t_b_96=249.848ns
.PARAM t_b_97=251.666667ns
.PARAM t_b_98=254.849ns
.PARAM t_b_99=256.666667ns
.PARAM t_b_100=259.85ns
.PARAM t_b_101=261.666667ns
.PARAM t_b_102=264.851ns
.PARAM t_b_103=266.666667ns
.PARAM t_b_104=269.852ns
.PARAM t_b_105=271.666667ns
.PARAM t_b_106=274.853ns
.PARAM t_b_107=276.666667ns
.PARAM t_b_108=279.854ns
.PARAM t_b_109=281.666667ns
.PARAM t_b_110=284.855ns
.PARAM t_b_111=286.666667ns
.PARAM t_b_112=289.856ns
.PARAM t_b_113=291.666667ns
.PARAM t_b_114=294.857ns
.PARAM t_b_115=296.666667ns
.PARAM t_b_116=299.858ns
.PARAM t_b_117=301.666667ns
.PARAM t_b_118=304.859ns
.PARAM t_b_119=306.666667ns
.PARAM t_b_120=309.86ns
.PARAM t_b_121=311.666667ns
.PARAM t_b_122=314.861ns
.PARAM t_b_123=316.666667ns
.PARAM t_b_124=319.862ns
.PARAM t_b_125=321.666667ns
.PARAM t_b_126=324.863ns
.PARAM t_b_127=326.666667ns
.PARAM t_b_128=329.864ns
.PARAM t_b_129=331.666667ns
.PARAM t_b_130=334.865ns
.PARAM t_b_131=336.666667ns
.PARAM t_b_132=339.866ns
.PARAM t_b_133=341.666667ns
.PARAM t_b_134=344.867ns
.PARAM t_b_135=346.666667ns
.PARAM t_b_136=349.868ns
.PARAM t_b_137=351.666667ns
.PARAM t_b_138=354.869ns
.PARAM t_b_139=356.666667ns
.PARAM t_b_140=359.87ns
.PARAM t_b_141=361.666667ns
.PARAM t_b_142=364.871ns
.PARAM t_b_143=366.666667ns
.PARAM t_b_144=369.872ns
.PARAM t_b_145=371.666667ns
.PARAM t_b_146=374.873ns
.PARAM t_b_147=376.666667ns
.PARAM t_b_148=379.874ns
.PARAM t_b_149=381.666667ns
.PARAM t_b_150=384.875ns
.PARAM t_b_151=386.666667ns
.PARAM t_b_152=389.876ns
.PARAM t_b_153=391.666667ns
.PARAM t_b_154=394.877ns
.PARAM t_b_155=396.666667ns
.PARAM t_b_156=399.878ns
.PARAM t_b_157=401.666667ns
.PARAM t_b_158=404.879ns
.PARAM t_b_159=406.666667ns
.PARAM t_b_160=409.88ns
.PARAM t_b_161=411.666667ns
.PARAM t_b_162=414.881ns
.PARAM t_b_163=416.666667ns
.PARAM t_b_164=419.882ns
.PARAM t_b_165=421.666667ns
.PARAM t_b_166=424.883ns
.PARAM t_b_167=426.666667ns
.PARAM t_b_168=429.884ns
.PARAM t_b_169=431.666667ns
.PARAM t_b_170=434.885ns
.PARAM t_b_171=436.666667ns
.PARAM t_b_172=439.886ns
.PARAM t_b_173=441.666667ns
.PARAM t_b_174=444.887ns
.PARAM t_b_175=446.666667ns
.PARAM t_b_176=449.888ns
.PARAM t_b_177=451.666667ns
.PARAM t_b_178=454.889ns
.PARAM t_b_179=456.666667ns
.PARAM t_b_180=459.89ns
.PARAM t_b_181=461.666667ns
.PARAM t_b_182=464.891ns
.PARAM t_b_183=466.666667ns
.PARAM t_b_184=469.892ns
.PARAM t_b_185=471.666667ns
.PARAM t_b_186=474.893ns
.PARAM t_b_187=476.666667ns
.PARAM t_b_188=479.894ns
.PARAM t_b_189=481.666667ns
.PARAM t_b_190=484.895ns
.PARAM t_b_191=486.666667ns
.PARAM t_b_192=489.896ns
.PARAM t_b_193=491.666667ns
.PARAM t_b_194=494.897ns
.PARAM t_b_195=496.666667ns
.PARAM t_b_196=499.898ns
.PARAM t_b_197=501.666667ns
.PARAM t_b_198=504.899ns
.PARAM t_b_199=506.666667ns
.PARAM t_b_200=509.9ns
.PARAM t_b_201=511.666667ns
.PARAM t_b_202=514.901ns
.PARAM t_b_203=516.666667ns
.PARAM t_b_204=519.902ns
.PARAM t_b_205=521.666667ns
.PARAM t_b_206=524.903ns
.PARAM t_b_207=526.666667ns
.PARAM t_b_208=529.904ns
.PARAM t_b_209=531.666667ns
.PARAM t_b_210=534.905ns
.PARAM t_b_211=536.666667ns
.PARAM t_b_212=539.906ns
.PARAM t_b_213=541.666667ns
.PARAM t_b_214=544.907ns
.PARAM t_b_215=546.666667ns
.PARAM t_b_216=549.908ns
.PARAM t_b_217=551.666667ns
.PARAM t_b_218=554.909ns
.PARAM t_b_219=556.666667ns
.PARAM t_b_220=559.91ns
.PARAM t_b_221=561.666667ns
.PARAM t_b_222=564.911ns
.PARAM t_b_223=566.666667ns
.PARAM t_b_224=569.912ns
.PARAM t_b_225=571.666667ns
.PARAM t_b_226=574.913ns
.PARAM t_b_227=576.666667ns
.PARAM t_b_228=579.914ns
.PARAM t_b_229=581.666667ns
.PARAM t_b_230=584.915ns
.PARAM t_b_231=586.666667ns
.PARAM t_b_232=589.916ns
.PARAM t_b_233=591.666667ns
.PARAM t_b_234=594.917ns
.PARAM t_b_235=596.666667ns
.PARAM t_b_236=599.918ns
.PARAM t_b_237=601.666667ns
.PARAM t_b_238=604.919ns
.PARAM t_b_239=606.666667ns
.PARAM t_b_240=609.92ns
.PARAM t_b_241=611.666667ns
.PARAM t_b_242=614.921ns
.PARAM t_b_243=616.666667ns
.PARAM t_b_244=619.922ns
.PARAM t_b_245=621.666667ns
.PARAM t_b_246=624.923ns
.PARAM t_b_247=626.666667ns
.PARAM t_b_248=629.924ns
.PARAM t_b_249=631.666667ns
.PARAM t_b_250=634.925ns
.PARAM t_b_251=636.666667ns
.PARAM t_b_252=639.926ns
.PARAM t_b_253=641.666667ns
.PARAM t_b_254=644.927ns
.PARAM t_b_255=646.666667ns
.PARAM t_b_256=649.928ns
.PARAM t_b_257=651.666667ns
.PARAM t_b_258=654.929ns
.PARAM t_b_259=656.666667ns
.PARAM t_b_260=659.93ns
.PARAM t_b_261=661.666667ns
.PARAM t_b_262=664.931ns
.PARAM t_b_263=666.666667ns
.PARAM t_b_264=669.932ns
.PARAM t_b_265=671.666667ns
.PARAM t_b_266=674.933ns
.PARAM t_b_267=676.666667ns
.PARAM t_b_268=679.934ns
.PARAM t_b_269=681.666667ns
.PARAM t_b_270=684.935ns
.PARAM t_b_271=686.666667ns
.PARAM t_b_272=689.936ns
.PARAM t_b_273=691.666667ns
.PARAM t_b_274=694.937ns
.PARAM t_b_275=696.666667ns
.PARAM t_b_276=699.938ns
.PARAM t_b_277=701.666667ns
.PARAM t_b_278=704.939ns
.PARAM t_b_279=706.666667ns
.PARAM t_b_280=709.94ns
.PARAM t_b_281=711.666667ns
.PARAM t_b_282=714.941ns
.PARAM t_b_283=716.666667ns
.PARAM t_b_284=719.942ns
.PARAM t_b_285=721.666667ns
.PARAM t_b_286=724.943ns
.PARAM t_b_287=726.666667ns
.PARAM t_b_288=729.944ns
.PARAM t_b_289=731.666667ns
.PARAM t_b_290=734.945ns
.PARAM t_b_291=736.666667ns
.PARAM t_b_292=739.946ns
.PARAM t_b_293=741.666667ns
.PARAM t_b_294=744.947ns
.PARAM t_b_295=746.666667ns
.PARAM t_b_296=749.948ns
.PARAM t_b_297=751.666667ns
.PARAM t_b_298=754.949ns
.PARAM t_b_299=756.666667ns
.PARAM t_b_300=759.95ns
.PARAM t_b_301=761.666667ns
.PARAM t_b_302=764.951ns
.PARAM t_b_303=766.666667ns
.PARAM t_b_304=769.952ns
.PARAM t_b_305=771.666667ns
.PARAM t_b_306=774.953ns
.PARAM t_b_307=776.666667ns
.PARAM t_b_308=779.954ns
.PARAM t_b_309=781.666667ns
.PARAM t_b_310=784.955ns
.PARAM t_b_311=786.666667ns
.PARAM t_b_312=789.956ns
.PARAM t_b_313=791.666667ns
.PARAM t_b_314=794.957ns
.PARAM t_b_315=796.666667ns
.PARAM t_b_316=799.958ns
.PARAM t_b_317=801.666667ns
.PARAM t_b_318=804.959ns
.PARAM t_b_319=806.666667ns
.PARAM t_b_320=809.96ns
.PARAM t_b_321=811.666667ns
.PARAM t_b_322=814.961ns
.PARAM t_b_323=816.666667ns
.PARAM t_b_324=819.962ns
.PARAM t_b_325=821.666667ns
.PARAM t_b_326=824.963ns
.PARAM t_b_327=826.666667ns
.PARAM t_b_328=829.964ns
.PARAM t_b_329=831.666667ns
.PARAM t_b_330=834.965ns
.PARAM t_b_331=836.666667ns
.PARAM t_b_332=839.966ns
.PARAM t_b_333=841.666667ns
.PARAM t_b_334=844.967ns
.PARAM t_b_335=846.666667ns
.PARAM t_b_336=849.968ns
.PARAM t_b_337=851.666667ns
.PARAM t_b_338=854.969ns
.PARAM t_b_339=856.666667ns
.PARAM t_b_340=859.97ns
.PARAM t_b_341=861.666667ns
.PARAM t_b_342=864.971ns
.PARAM t_b_343=866.666667ns
.PARAM t_b_344=869.972ns
.PARAM t_b_345=871.666667ns
.PARAM t_b_346=874.973ns
.PARAM t_b_347=876.666667ns
.PARAM t_b_348=879.974ns
.PARAM t_b_349=881.666667ns
.PARAM t_b_350=884.975ns
.PARAM t_b_351=886.666667ns
.PARAM t_b_352=889.976ns
.PARAM t_b_353=891.666667ns
.PARAM t_b_354=894.977ns
.PARAM t_b_355=896.666667ns
.PARAM t_b_356=899.978ns
.PARAM t_b_357=901.666667ns
.PARAM t_b_358=904.979ns
.PARAM t_b_359=906.666667ns
.PARAM t_b_360=909.98ns
.PARAM t_b_361=911.666667ns
.PARAM t_b_362=914.981ns
.PARAM t_b_363=916.666667ns
.PARAM t_b_364=919.982ns
.PARAM t_b_365=921.666667ns
.PARAM t_b_366=924.983ns
.PARAM t_b_367=926.666667ns
.PARAM t_b_368=929.984ns
.PARAM t_b_369=931.666667ns
.PARAM t_b_370=934.985ns
.PARAM t_b_371=936.666667ns
.PARAM t_b_372=939.986ns
.PARAM t_b_373=941.666667ns
.PARAM t_b_374=944.987ns
.PARAM t_b_375=946.666667ns
.PARAM t_b_376=949.988ns
.PARAM t_b_377=951.666667ns
.PARAM t_b_378=954.989ns
.PARAM t_b_379=956.666667ns
.PARAM t_b_380=959.99ns
.PARAM t_b_381=961.666667ns
.PARAM t_b_382=964.991ns
.PARAM t_b_383=966.666667ns
.PARAM t_b_384=969.992ns
.PARAM t_b_385=971.666667ns
.PARAM t_b_386=974.993ns
.PARAM t_b_387=976.666667ns
.PARAM t_b_388=979.994ns
.PARAM t_b_389=981.666667ns
.PARAM t_b_390=984.995ns
.PARAM t_b_391=986.666667ns
.PARAM t_b_392=989.996ns
.PARAM t_b_393=991.666667ns
.PARAM t_b_394=994.997ns
.PARAM t_b_395=996.666667ns
.PARAM t_b_396=999.998ns
.PARAM t_b_397=1001.666667ns
.PARAM t_b_398=1004.999ns
.PARAM t_b_399=1006.666667ns
.PARAM t_b_400=1010.0ns
.PARAM t_b_401=1011.666667ns
.PARAM t_b_402=1015.001ns
.PARAM t_b_403=1016.666667ns
.PARAM t_b_404=1020.002ns
.PARAM t_b_405=1021.666667ns
.PARAM t_b_406=1025.003ns
.PARAM t_b_407=1026.666667ns
.PARAM t_b_408=1030.004ns
.PARAM t_b_409=1031.666667ns
.PARAM t_b_410=1035.005ns
.PARAM t_b_411=1036.666667ns
.PARAM t_b_412=1040.006ns
.PARAM t_b_413=1041.666667ns
.PARAM t_b_414=1045.007ns
.PARAM t_b_415=1046.666667ns
.PARAM t_b_416=1050.008ns
.PARAM t_b_417=1051.666667ns
.PARAM t_b_418=1055.009ns
.PARAM t_b_419=1056.666667ns
.PARAM t_b_420=1060.01ns
.PARAM t_b_421=1061.666667ns
.PARAM t_b_422=1065.011ns
.PARAM t_b_423=1066.666667ns
.PARAM t_b_424=1070.012ns
.PARAM t_b_425=1071.666667ns
.PARAM t_b_426=1075.013ns
.PARAM t_b_427=1076.666667ns
.PARAM t_b_428=1080.014ns
.PARAM t_b_429=1081.666667ns
.PARAM t_b_430=1085.015ns
.PARAM t_b_431=1086.666667ns
.PARAM t_b_432=1090.016ns
.PARAM t_b_433=1091.666667ns
.PARAM t_b_434=1095.017ns
.PARAM t_b_435=1096.666667ns
.PARAM t_b_436=1100.018ns
.PARAM t_b_437=1101.666667ns
.PARAM t_b_438=1105.019ns
.PARAM t_b_439=1106.666667ns
.PARAM t_b_440=1110.02ns
.PARAM t_b_441=1111.666667ns
.PARAM t_b_442=1115.021ns
.PARAM t_b_443=1116.666667ns
.PARAM t_b_444=1120.022ns
.PARAM t_b_445=1121.666667ns
.PARAM t_b_446=1125.023ns
.PARAM t_b_447=1126.666667ns
.PARAM t_b_448=1130.024ns
.PARAM t_b_449=1131.666667ns
.PARAM t_b_450=1135.025ns
.PARAM t_b_451=1136.666667ns
.PARAM t_b_452=1140.026ns
.PARAM t_b_453=1141.666667ns
.PARAM t_b_454=1145.027ns
.PARAM t_b_455=1146.666667ns
.PARAM t_b_456=1150.028ns
.PARAM t_b_457=1151.666667ns
.PARAM t_b_458=1155.029ns
.PARAM t_b_459=1156.666667ns
.PARAM t_b_460=1160.03ns
.PARAM t_b_461=1161.666667ns
.PARAM t_b_462=1165.031ns
.PARAM t_b_463=1166.666667ns
.PARAM t_b_464=1170.032ns
.PARAM t_b_465=1171.666667ns
.PARAM t_b_466=1175.033ns
.PARAM t_b_467=1176.666667ns
.PARAM t_b_468=1180.034ns
.PARAM t_b_469=1181.666667ns
.PARAM t_b_470=1185.035ns
.PARAM t_b_471=1186.666667ns
.PARAM t_b_472=1190.036ns
.PARAM t_b_473=1191.666667ns
.PARAM t_b_474=1195.037ns
.PARAM t_b_475=1196.666667ns
.PARAM t_b_476=1200.038ns
.PARAM t_b_477=1201.666667ns
.PARAM t_b_478=1205.039ns
.PARAM t_b_479=1206.666667ns
.PARAM t_b_480=1210.04ns
.PARAM t_b_481=1211.666667ns
.PARAM t_b_482=1215.041ns
.PARAM t_b_483=1216.666667ns
.PARAM t_b_484=1220.042ns
.PARAM t_b_485=1221.666667ns
.PARAM t_b_486=1225.043ns
.PARAM t_b_487=1226.666667ns
.PARAM t_b_488=1230.044ns
.PARAM t_b_489=1231.666667ns
.PARAM t_b_490=1235.045ns
.PARAM t_b_491=1236.666667ns
.PARAM t_b_492=1240.046ns
.PARAM t_b_493=1241.666667ns
.PARAM t_b_494=1245.047ns
.PARAM t_b_495=1246.666667ns
.PARAM t_b_496=1250.048ns
.PARAM t_b_497=1251.666667ns
.PARAM t_b_498=1255.049ns
.PARAM t_b_499=1256.666667ns
.PARAM t_b_500=1260.05ns
.PARAM t_b_501=1261.666667ns
.PARAM t_b_502=1265.051ns
.PARAM t_b_503=1266.666667ns
.PARAM t_b_504=1270.052ns
.PARAM t_b_505=1271.666667ns
.PARAM t_b_506=1275.053ns
.PARAM t_b_507=1276.666667ns
.PARAM t_b_508=1280.054ns
.PARAM t_b_509=1281.666667ns
.PARAM t_b_510=1285.055ns
.PARAM t_b_511=1286.666667ns
.PARAM t_b_512=1290.056ns
.PARAM t_b_513=1291.666667ns
.PARAM t_b_514=1295.057ns
.PARAM t_b_515=1296.666667ns
.PARAM t_b_516=1300.058ns
.PARAM t_b_517=1301.666667ns
.PARAM t_b_518=1305.059ns
.PARAM t_b_519=1306.666667ns
.PARAM t_b_520=1310.06ns
.PARAM t_b_521=1311.666667ns
.PARAM t_b_522=1315.061ns
.PARAM t_b_523=1316.666667ns
.PARAM t_b_524=1320.062ns
.PARAM t_b_525=1321.666667ns
.PARAM t_b_526=1325.063ns
.PARAM t_b_527=1326.666667ns
.PARAM t_b_528=1330.064ns
.PARAM t_b_529=1331.666667ns
.PARAM t_b_530=1335.065ns
.PARAM t_b_531=1336.666667ns
.PARAM t_b_532=1340.066ns
.PARAM t_b_533=1341.666667ns
.PARAM t_b_534=1345.067ns
.PARAM t_b_535=1346.666667ns
.PARAM t_b_536=1350.068ns
.PARAM t_b_537=1351.666667ns
.PARAM t_b_538=1355.069ns
.PARAM t_b_539=1356.666667ns
.PARAM t_b_540=1360.07ns
.PARAM t_b_541=1361.666667ns
.PARAM t_b_542=1365.071ns
.PARAM t_b_543=1366.666667ns
.PARAM t_b_544=1370.072ns
.PARAM t_b_545=1371.666667ns
.PARAM t_b_546=1375.073ns
.PARAM t_b_547=1376.666667ns
.PARAM t_b_548=1380.074ns
.PARAM t_b_549=1381.666667ns
.PARAM t_b_550=1385.075ns
.PARAM t_b_551=1386.666667ns
.PARAM t_b_552=1390.076ns
.PARAM t_b_553=1391.666667ns
.PARAM t_b_554=1395.077ns
.PARAM t_b_555=1396.666667ns
.PARAM t_b_556=1400.078ns
.PARAM t_b_557=1401.666667ns
.PARAM t_b_558=1405.079ns
.PARAM t_b_559=1406.666667ns
.PARAM t_b_560=1410.08ns
.PARAM t_b_561=1411.666667ns
.PARAM t_b_562=1415.081ns
.PARAM t_b_563=1416.666667ns
.PARAM t_b_564=1420.082ns
.PARAM t_b_565=1421.666667ns
.PARAM t_b_566=1425.083ns
.PARAM t_b_567=1426.666667ns
.PARAM t_b_568=1430.084ns
.PARAM t_b_569=1431.666667ns
.PARAM t_b_570=1435.085ns
.PARAM t_b_571=1436.666667ns
.PARAM t_b_572=1440.086ns
.PARAM t_b_573=1441.666667ns
.PARAM t_b_574=1445.087ns
.PARAM t_b_575=1446.666667ns
.PARAM t_b_576=1450.088ns
.PARAM t_b_577=1451.666667ns
.PARAM t_b_578=1455.089ns
.PARAM t_b_579=1456.666667ns
.PARAM t_b_580=1460.09ns
.PARAM t_b_581=1461.666667ns
.PARAM t_b_582=1465.091ns
.PARAM t_b_583=1466.666667ns
.PARAM t_b_584=1470.092ns
.PARAM t_b_585=1471.666667ns
.PARAM t_b_586=1475.093ns
.PARAM t_b_587=1476.666667ns
.PARAM t_b_588=1480.094ns
.PARAM t_b_589=1481.666667ns
.PARAM t_b_590=1485.095ns
.PARAM t_b_591=1486.666667ns
.PARAM t_b_592=1490.096ns
.PARAM t_b_593=1491.666667ns
.PARAM t_b_594=1495.097ns
.PARAM t_b_595=1496.666667ns
.PARAM t_b_596=1500.098ns
.PARAM t_b_597=1501.666667ns
.PARAM t_b_598=1505.099ns
.PARAM t_b_599=1506.666667ns
.PARAM t_b_600=1510.1ns
.PARAM t_b_601=1511.666667ns
.PARAM t_b_602=1515.101ns
.PARAM t_b_603=1516.666667ns
.PARAM t_b_604=1520.102ns
.PARAM t_b_605=1521.666667ns
.PARAM t_b_606=1525.103ns
.PARAM t_b_607=1526.666667ns
.PARAM t_b_608=1530.104ns
.PARAM t_b_609=1531.666667ns
.PARAM t_b_610=1535.105ns
.PARAM t_b_611=1536.666667ns
.PARAM t_b_612=1540.106ns
.PARAM t_b_613=1541.666667ns
.PARAM t_b_614=1545.107ns
.PARAM t_b_615=1546.666667ns
.PARAM t_b_616=1550.108ns
.PARAM t_b_617=1551.666667ns
.PARAM t_b_618=1555.109ns
.PARAM t_b_619=1556.666667ns
.PARAM t_b_620=1560.11ns
.PARAM t_b_621=1561.666667ns
.PARAM t_b_622=1565.111ns
.PARAM t_b_623=1566.666667ns
.PARAM t_b_624=1570.112ns
.PARAM t_b_625=1571.666667ns
.PARAM t_b_626=1575.113ns
.PARAM t_b_627=1576.666667ns
.PARAM t_b_628=1580.114ns
.PARAM t_b_629=1581.666667ns
.PARAM t_b_630=1585.115ns
.PARAM t_b_631=1586.666667ns
.PARAM t_b_632=1590.116ns
.PARAM t_b_633=1591.666667ns
.PARAM t_b_634=1595.117ns
.PARAM t_b_635=1596.666667ns
.PARAM t_b_636=1600.118ns
.PARAM t_b_637=1601.666667ns
.PARAM t_b_638=1605.119ns
.PARAM t_b_639=1606.666667ns
.PARAM t_b_640=1610.12ns
.PARAM t_b_641=1611.666667ns
.PARAM t_b_642=1615.121ns
.PARAM t_b_643=1616.666667ns
.PARAM t_b_644=1620.122ns
.PARAM t_b_645=1621.666667ns
.PARAM t_b_646=1625.123ns
.PARAM t_b_647=1626.666667ns
.PARAM t_b_648=1630.124ns
.PARAM t_b_649=1631.666667ns
.PARAM t_b_650=1635.125ns
.PARAM t_b_651=1636.666667ns
.PARAM t_b_652=1640.126ns
.PARAM t_b_653=1641.666667ns
.PARAM t_b_654=1645.127ns
.PARAM t_b_655=1646.666667ns
.PARAM t_b_656=1650.128ns
.PARAM t_b_657=1651.666667ns
.PARAM t_b_658=1655.129ns
.PARAM t_b_659=1656.666667ns
.PARAM t_b_660=1660.13ns
.PARAM t_b_661=1661.666667ns
.PARAM t_b_662=1665.131ns
.PARAM t_b_663=1666.666667ns
.PARAM t_b_664=1670.132ns
.PARAM t_b_665=1671.666667ns
.PARAM t_b_666=1675.133ns
.PARAM t_b_667=1676.666667ns
.PARAM t_b_668=1680.134ns
.PARAM t_b_669=1681.666667ns
.PARAM t_b_670=1685.135ns
.PARAM t_b_671=1686.666667ns
.PARAM t_b_672=1690.136ns
.PARAM t_b_673=1691.666667ns
.PARAM t_b_674=1695.137ns
.PARAM t_b_675=1696.666667ns
.PARAM t_b_676=1700.138ns
.PARAM t_b_677=1701.666667ns
.PARAM t_b_678=1705.139ns
.PARAM t_b_679=1706.666667ns
.PARAM t_b_680=1710.14ns
.PARAM t_b_681=1711.666667ns
.PARAM t_b_682=1715.141ns
.PARAM t_b_683=1716.666667ns
.PARAM t_b_684=1720.142ns
.PARAM t_b_685=1721.666667ns
.PARAM t_b_686=1725.143ns
.PARAM t_b_687=1726.666667ns
.PARAM t_b_688=1730.144ns
.PARAM t_b_689=1731.666667ns
.PARAM t_b_690=1735.145ns
.PARAM t_b_691=1736.666667ns
.PARAM t_b_692=1740.146ns
.PARAM t_b_693=1741.666667ns
.PARAM t_b_694=1745.147ns
.PARAM t_b_695=1746.666667ns
.PARAM t_b_696=1750.148ns
.PARAM t_b_697=1751.666667ns
.PARAM t_b_698=1755.149ns
.PARAM t_b_699=1756.666667ns
.PARAM t_b_700=1760.15ns
.PARAM t_b_701=1761.666667ns
.PARAM t_b_702=1765.151ns
.PARAM t_b_703=1766.666667ns
.PARAM t_b_704=1770.152ns
.PARAM t_b_705=1771.666667ns
.PARAM t_b_706=1775.153ns
.PARAM t_b_707=1776.666667ns
.PARAM t_b_708=1780.154ns
.PARAM t_b_709=1781.666667ns
.PARAM t_b_710=1785.155ns
.PARAM t_b_711=1786.666667ns
.PARAM t_b_712=1790.156ns
.PARAM t_b_713=1791.666667ns
.PARAM t_b_714=1795.157ns
.PARAM t_b_715=1796.666667ns
.PARAM t_b_716=1800.158ns
.PARAM t_b_717=1801.666667ns
.PARAM t_b_718=1805.159ns
.PARAM t_b_719=1806.666667ns
.PARAM t_b_720=1810.16ns
.PARAM t_b_721=1811.666667ns
.PARAM t_b_722=1815.161ns
.PARAM t_b_723=1816.666667ns
.PARAM t_b_724=1820.162ns
.PARAM t_b_725=1821.666667ns
.PARAM t_b_726=1825.163ns
.PARAM t_b_727=1826.666667ns
.PARAM t_b_728=1830.164ns
.PARAM t_b_729=1831.666667ns
.PARAM t_b_730=1835.165ns
.PARAM t_b_731=1836.666667ns
.PARAM t_b_732=1840.166ns
.PARAM t_b_733=1841.666667ns
.PARAM t_b_734=1845.167ns
.PARAM t_b_735=1846.666667ns
.PARAM t_b_736=1850.168ns
.PARAM t_b_737=1851.666667ns
.PARAM t_b_738=1855.169ns
.PARAM t_b_739=1856.666667ns
.PARAM t_b_740=1860.17ns
.PARAM t_b_741=1861.666667ns
.PARAM t_b_742=1865.171ns
.PARAM t_b_743=1866.666667ns
.PARAM t_b_744=1870.172ns
.PARAM t_b_745=1871.666667ns
.PARAM t_b_746=1875.173ns
.PARAM t_b_747=1876.666667ns
.PARAM t_b_748=1880.174ns
.PARAM t_b_749=1881.666667ns
.PARAM t_b_750=1885.175ns
.PARAM t_b_751=1886.666667ns
.PARAM t_b_752=1890.176ns
.PARAM t_b_753=1891.666667ns
.PARAM t_b_754=1895.177ns
.PARAM t_b_755=1896.666667ns
.PARAM t_b_756=1900.178ns
.PARAM t_b_757=1901.666667ns
.PARAM t_b_758=1905.179ns
.PARAM t_b_759=1906.666667ns
.PARAM t_b_760=1910.18ns
.PARAM t_b_761=1911.666667ns
.PARAM t_b_762=1915.181ns
.PARAM t_b_763=1916.666667ns
.PARAM t_b_764=1920.182ns
.PARAM t_b_765=1921.666667ns
.PARAM t_b_766=1925.183ns
.PARAM t_b_767=1926.666667ns
.PARAM t_b_768=1930.184ns
.PARAM t_b_769=1931.666667ns
.PARAM t_b_770=1935.185ns
.PARAM t_b_771=1936.666667ns
.PARAM t_b_772=1940.186ns
.PARAM t_b_773=1941.666667ns
.PARAM t_b_774=1945.187ns
.PARAM t_b_775=1946.666667ns
.PARAM t_b_776=1950.188ns
.PARAM t_b_777=1951.666667ns
.PARAM t_b_778=1955.189ns
.PARAM t_b_779=1956.666667ns
.PARAM t_b_780=1960.19ns
.PARAM t_b_781=1961.666667ns
.PARAM t_b_782=1965.191ns
.PARAM t_b_783=1966.666667ns
.PARAM t_b_784=1970.192ns
.PARAM t_b_785=1971.666667ns
.PARAM t_b_786=1975.193ns
.PARAM t_b_787=1976.666667ns
.PARAM t_b_788=1980.194ns
.PARAM t_b_789=1981.666667ns
.PARAM t_b_790=1985.195ns
.PARAM t_b_791=1986.666667ns
.PARAM t_b_792=1990.196ns
.PARAM t_b_793=1991.666667ns
.PARAM t_b_794=1995.197ns
.PARAM t_b_795=1996.666667ns
.PARAM t_b_796=2000.198ns
.PARAM t_b_797=2001.666667ns
.PARAM t_b_798=2005.199ns
.PARAM t_b_799=2006.666667ns



VINA Input_A GND PWL 0ns baseVal t_init0 baseVal 't_init0+slope' peakVal t_init1 peakVal 't_init1+slope' baseVal
+ t_a_0 peakVal 't_a_0+slope' baseVal
+ t_a_1 baseVal 't_a_1+slope' peakVal
+ t_a_2 peakVal 't_a_2+slope' baseVal
+ t_a_3 baseVal 't_a_3+slope' peakVal
+ t_a_4 peakVal 't_a_4+slope' baseVal
+ t_a_5 baseVal 't_a_5+slope' peakVal
+ t_a_6 peakVal 't_a_6+slope' baseVal
+ t_a_7 baseVal 't_a_7+slope' peakVal
+ t_a_8 peakVal 't_a_8+slope' baseVal
+ t_a_9 baseVal 't_a_9+slope' peakVal
+ t_a_10 peakVal 't_a_10+slope' baseVal
+ t_a_11 baseVal 't_a_11+slope' peakVal
+ t_a_12 peakVal 't_a_12+slope' baseVal
+ t_a_13 baseVal 't_a_13+slope' peakVal
+ t_a_14 peakVal 't_a_14+slope' baseVal
+ t_a_15 baseVal 't_a_15+slope' peakVal
+ t_a_16 peakVal 't_a_16+slope' baseVal
+ t_a_17 baseVal 't_a_17+slope' peakVal
+ t_a_18 peakVal 't_a_18+slope' baseVal
+ t_a_19 baseVal 't_a_19+slope' peakVal
+ t_a_20 peakVal 't_a_20+slope' baseVal
+ t_a_21 baseVal 't_a_21+slope' peakVal
+ t_a_22 peakVal 't_a_22+slope' baseVal
+ t_a_23 baseVal 't_a_23+slope' peakVal
+ t_a_24 peakVal 't_a_24+slope' baseVal
+ t_a_25 baseVal 't_a_25+slope' peakVal
+ t_a_26 peakVal 't_a_26+slope' baseVal
+ t_a_27 baseVal 't_a_27+slope' peakVal
+ t_a_28 peakVal 't_a_28+slope' baseVal
+ t_a_29 baseVal 't_a_29+slope' peakVal
+ t_a_30 peakVal 't_a_30+slope' baseVal
+ t_a_31 baseVal 't_a_31+slope' peakVal
+ t_a_32 peakVal 't_a_32+slope' baseVal
+ t_a_33 baseVal 't_a_33+slope' peakVal
+ t_a_34 peakVal 't_a_34+slope' baseVal
+ t_a_35 baseVal 't_a_35+slope' peakVal
+ t_a_36 peakVal 't_a_36+slope' baseVal
+ t_a_37 baseVal 't_a_37+slope' peakVal
+ t_a_38 peakVal 't_a_38+slope' baseVal
+ t_a_39 baseVal 't_a_39+slope' peakVal
+ t_a_40 peakVal 't_a_40+slope' baseVal
+ t_a_41 baseVal 't_a_41+slope' peakVal
+ t_a_42 peakVal 't_a_42+slope' baseVal
+ t_a_43 baseVal 't_a_43+slope' peakVal
+ t_a_44 peakVal 't_a_44+slope' baseVal
+ t_a_45 baseVal 't_a_45+slope' peakVal
+ t_a_46 peakVal 't_a_46+slope' baseVal
+ t_a_47 baseVal 't_a_47+slope' peakVal
+ t_a_48 peakVal 't_a_48+slope' baseVal
+ t_a_49 baseVal 't_a_49+slope' peakVal
+ t_a_50 peakVal 't_a_50+slope' baseVal
+ t_a_51 baseVal 't_a_51+slope' peakVal
+ t_a_52 peakVal 't_a_52+slope' baseVal
+ t_a_53 baseVal 't_a_53+slope' peakVal
+ t_a_54 peakVal 't_a_54+slope' baseVal
+ t_a_55 baseVal 't_a_55+slope' peakVal
+ t_a_56 peakVal 't_a_56+slope' baseVal
+ t_a_57 baseVal 't_a_57+slope' peakVal
+ t_a_58 peakVal 't_a_58+slope' baseVal
+ t_a_59 baseVal 't_a_59+slope' peakVal
+ t_a_60 peakVal 't_a_60+slope' baseVal
+ t_a_61 baseVal 't_a_61+slope' peakVal
+ t_a_62 peakVal 't_a_62+slope' baseVal
+ t_a_63 baseVal 't_a_63+slope' peakVal
+ t_a_64 peakVal 't_a_64+slope' baseVal
+ t_a_65 baseVal 't_a_65+slope' peakVal
+ t_a_66 peakVal 't_a_66+slope' baseVal
+ t_a_67 baseVal 't_a_67+slope' peakVal
+ t_a_68 peakVal 't_a_68+slope' baseVal
+ t_a_69 baseVal 't_a_69+slope' peakVal
+ t_a_70 peakVal 't_a_70+slope' baseVal
+ t_a_71 baseVal 't_a_71+slope' peakVal
+ t_a_72 peakVal 't_a_72+slope' baseVal
+ t_a_73 baseVal 't_a_73+slope' peakVal
+ t_a_74 peakVal 't_a_74+slope' baseVal
+ t_a_75 baseVal 't_a_75+slope' peakVal
+ t_a_76 peakVal 't_a_76+slope' baseVal
+ t_a_77 baseVal 't_a_77+slope' peakVal
+ t_a_78 peakVal 't_a_78+slope' baseVal
+ t_a_79 baseVal 't_a_79+slope' peakVal
+ t_a_80 peakVal 't_a_80+slope' baseVal
+ t_a_81 baseVal 't_a_81+slope' peakVal
+ t_a_82 peakVal 't_a_82+slope' baseVal
+ t_a_83 baseVal 't_a_83+slope' peakVal
+ t_a_84 peakVal 't_a_84+slope' baseVal
+ t_a_85 baseVal 't_a_85+slope' peakVal
+ t_a_86 peakVal 't_a_86+slope' baseVal
+ t_a_87 baseVal 't_a_87+slope' peakVal
+ t_a_88 peakVal 't_a_88+slope' baseVal
+ t_a_89 baseVal 't_a_89+slope' peakVal
+ t_a_90 peakVal 't_a_90+slope' baseVal
+ t_a_91 baseVal 't_a_91+slope' peakVal
+ t_a_92 peakVal 't_a_92+slope' baseVal
+ t_a_93 baseVal 't_a_93+slope' peakVal
+ t_a_94 peakVal 't_a_94+slope' baseVal
+ t_a_95 baseVal 't_a_95+slope' peakVal
+ t_a_96 peakVal 't_a_96+slope' baseVal
+ t_a_97 baseVal 't_a_97+slope' peakVal
+ t_a_98 peakVal 't_a_98+slope' baseVal
+ t_a_99 baseVal 't_a_99+slope' peakVal
+ t_a_100 peakVal 't_a_100+slope' baseVal
+ t_a_101 baseVal 't_a_101+slope' peakVal
+ t_a_102 peakVal 't_a_102+slope' baseVal
+ t_a_103 baseVal 't_a_103+slope' peakVal
+ t_a_104 peakVal 't_a_104+slope' baseVal
+ t_a_105 baseVal 't_a_105+slope' peakVal
+ t_a_106 peakVal 't_a_106+slope' baseVal
+ t_a_107 baseVal 't_a_107+slope' peakVal
+ t_a_108 peakVal 't_a_108+slope' baseVal
+ t_a_109 baseVal 't_a_109+slope' peakVal
+ t_a_110 peakVal 't_a_110+slope' baseVal
+ t_a_111 baseVal 't_a_111+slope' peakVal
+ t_a_112 peakVal 't_a_112+slope' baseVal
+ t_a_113 baseVal 't_a_113+slope' peakVal
+ t_a_114 peakVal 't_a_114+slope' baseVal
+ t_a_115 baseVal 't_a_115+slope' peakVal
+ t_a_116 peakVal 't_a_116+slope' baseVal
+ t_a_117 baseVal 't_a_117+slope' peakVal
+ t_a_118 peakVal 't_a_118+slope' baseVal
+ t_a_119 baseVal 't_a_119+slope' peakVal
+ t_a_120 peakVal 't_a_120+slope' baseVal
+ t_a_121 baseVal 't_a_121+slope' peakVal
+ t_a_122 peakVal 't_a_122+slope' baseVal
+ t_a_123 baseVal 't_a_123+slope' peakVal
+ t_a_124 peakVal 't_a_124+slope' baseVal
+ t_a_125 baseVal 't_a_125+slope' peakVal
+ t_a_126 peakVal 't_a_126+slope' baseVal
+ t_a_127 baseVal 't_a_127+slope' peakVal
+ t_a_128 peakVal 't_a_128+slope' baseVal
+ t_a_129 baseVal 't_a_129+slope' peakVal
+ t_a_130 peakVal 't_a_130+slope' baseVal
+ t_a_131 baseVal 't_a_131+slope' peakVal
+ t_a_132 peakVal 't_a_132+slope' baseVal
+ t_a_133 baseVal 't_a_133+slope' peakVal
+ t_a_134 peakVal 't_a_134+slope' baseVal
+ t_a_135 baseVal 't_a_135+slope' peakVal
+ t_a_136 peakVal 't_a_136+slope' baseVal
+ t_a_137 baseVal 't_a_137+slope' peakVal
+ t_a_138 peakVal 't_a_138+slope' baseVal
+ t_a_139 baseVal 't_a_139+slope' peakVal
+ t_a_140 peakVal 't_a_140+slope' baseVal
+ t_a_141 baseVal 't_a_141+slope' peakVal
+ t_a_142 peakVal 't_a_142+slope' baseVal
+ t_a_143 baseVal 't_a_143+slope' peakVal
+ t_a_144 peakVal 't_a_144+slope' baseVal
+ t_a_145 baseVal 't_a_145+slope' peakVal
+ t_a_146 peakVal 't_a_146+slope' baseVal
+ t_a_147 baseVal 't_a_147+slope' peakVal
+ t_a_148 peakVal 't_a_148+slope' baseVal
+ t_a_149 baseVal 't_a_149+slope' peakVal
+ t_a_150 peakVal 't_a_150+slope' baseVal
+ t_a_151 baseVal 't_a_151+slope' peakVal
+ t_a_152 peakVal 't_a_152+slope' baseVal
+ t_a_153 baseVal 't_a_153+slope' peakVal
+ t_a_154 peakVal 't_a_154+slope' baseVal
+ t_a_155 baseVal 't_a_155+slope' peakVal
+ t_a_156 peakVal 't_a_156+slope' baseVal
+ t_a_157 baseVal 't_a_157+slope' peakVal
+ t_a_158 peakVal 't_a_158+slope' baseVal
+ t_a_159 baseVal 't_a_159+slope' peakVal
+ t_a_160 peakVal 't_a_160+slope' baseVal
+ t_a_161 baseVal 't_a_161+slope' peakVal
+ t_a_162 peakVal 't_a_162+slope' baseVal
+ t_a_163 baseVal 't_a_163+slope' peakVal
+ t_a_164 peakVal 't_a_164+slope' baseVal
+ t_a_165 baseVal 't_a_165+slope' peakVal
+ t_a_166 peakVal 't_a_166+slope' baseVal
+ t_a_167 baseVal 't_a_167+slope' peakVal
+ t_a_168 peakVal 't_a_168+slope' baseVal
+ t_a_169 baseVal 't_a_169+slope' peakVal
+ t_a_170 peakVal 't_a_170+slope' baseVal
+ t_a_171 baseVal 't_a_171+slope' peakVal
+ t_a_172 peakVal 't_a_172+slope' baseVal
+ t_a_173 baseVal 't_a_173+slope' peakVal
+ t_a_174 peakVal 't_a_174+slope' baseVal
+ t_a_175 baseVal 't_a_175+slope' peakVal
+ t_a_176 peakVal 't_a_176+slope' baseVal
+ t_a_177 baseVal 't_a_177+slope' peakVal
+ t_a_178 peakVal 't_a_178+slope' baseVal
+ t_a_179 baseVal 't_a_179+slope' peakVal
+ t_a_180 peakVal 't_a_180+slope' baseVal
+ t_a_181 baseVal 't_a_181+slope' peakVal
+ t_a_182 peakVal 't_a_182+slope' baseVal
+ t_a_183 baseVal 't_a_183+slope' peakVal
+ t_a_184 peakVal 't_a_184+slope' baseVal
+ t_a_185 baseVal 't_a_185+slope' peakVal
+ t_a_186 peakVal 't_a_186+slope' baseVal
+ t_a_187 baseVal 't_a_187+slope' peakVal
+ t_a_188 peakVal 't_a_188+slope' baseVal
+ t_a_189 baseVal 't_a_189+slope' peakVal
+ t_a_190 peakVal 't_a_190+slope' baseVal
+ t_a_191 baseVal 't_a_191+slope' peakVal
+ t_a_192 peakVal 't_a_192+slope' baseVal
+ t_a_193 baseVal 't_a_193+slope' peakVal
+ t_a_194 peakVal 't_a_194+slope' baseVal
+ t_a_195 baseVal 't_a_195+slope' peakVal
+ t_a_196 peakVal 't_a_196+slope' baseVal
+ t_a_197 baseVal 't_a_197+slope' peakVal
+ t_a_198 peakVal 't_a_198+slope' baseVal
+ t_a_199 baseVal 't_a_199+slope' peakVal
+ t_a_200 peakVal 't_a_200+slope' baseVal
+ t_a_201 baseVal 't_a_201+slope' peakVal
+ t_a_202 peakVal 't_a_202+slope' baseVal
+ t_a_203 baseVal 't_a_203+slope' peakVal
+ t_a_204 peakVal 't_a_204+slope' baseVal
+ t_a_205 baseVal 't_a_205+slope' peakVal
+ t_a_206 peakVal 't_a_206+slope' baseVal
+ t_a_207 baseVal 't_a_207+slope' peakVal
+ t_a_208 peakVal 't_a_208+slope' baseVal
+ t_a_209 baseVal 't_a_209+slope' peakVal
+ t_a_210 peakVal 't_a_210+slope' baseVal
+ t_a_211 baseVal 't_a_211+slope' peakVal
+ t_a_212 peakVal 't_a_212+slope' baseVal
+ t_a_213 baseVal 't_a_213+slope' peakVal
+ t_a_214 peakVal 't_a_214+slope' baseVal
+ t_a_215 baseVal 't_a_215+slope' peakVal
+ t_a_216 peakVal 't_a_216+slope' baseVal
+ t_a_217 baseVal 't_a_217+slope' peakVal
+ t_a_218 peakVal 't_a_218+slope' baseVal
+ t_a_219 baseVal 't_a_219+slope' peakVal
+ t_a_220 peakVal 't_a_220+slope' baseVal
+ t_a_221 baseVal 't_a_221+slope' peakVal
+ t_a_222 peakVal 't_a_222+slope' baseVal
+ t_a_223 baseVal 't_a_223+slope' peakVal
+ t_a_224 peakVal 't_a_224+slope' baseVal
+ t_a_225 baseVal 't_a_225+slope' peakVal
+ t_a_226 peakVal 't_a_226+slope' baseVal
+ t_a_227 baseVal 't_a_227+slope' peakVal
+ t_a_228 peakVal 't_a_228+slope' baseVal
+ t_a_229 baseVal 't_a_229+slope' peakVal
+ t_a_230 peakVal 't_a_230+slope' baseVal
+ t_a_231 baseVal 't_a_231+slope' peakVal
+ t_a_232 peakVal 't_a_232+slope' baseVal
+ t_a_233 baseVal 't_a_233+slope' peakVal
+ t_a_234 peakVal 't_a_234+slope' baseVal
+ t_a_235 baseVal 't_a_235+slope' peakVal
+ t_a_236 peakVal 't_a_236+slope' baseVal
+ t_a_237 baseVal 't_a_237+slope' peakVal
+ t_a_238 peakVal 't_a_238+slope' baseVal
+ t_a_239 baseVal 't_a_239+slope' peakVal
+ t_a_240 peakVal 't_a_240+slope' baseVal
+ t_a_241 baseVal 't_a_241+slope' peakVal
+ t_a_242 peakVal 't_a_242+slope' baseVal
+ t_a_243 baseVal 't_a_243+slope' peakVal
+ t_a_244 peakVal 't_a_244+slope' baseVal
+ t_a_245 baseVal 't_a_245+slope' peakVal
+ t_a_246 peakVal 't_a_246+slope' baseVal
+ t_a_247 baseVal 't_a_247+slope' peakVal
+ t_a_248 peakVal 't_a_248+slope' baseVal
+ t_a_249 baseVal 't_a_249+slope' peakVal
+ t_a_250 peakVal 't_a_250+slope' baseVal
+ t_a_251 baseVal 't_a_251+slope' peakVal
+ t_a_252 peakVal 't_a_252+slope' baseVal
+ t_a_253 baseVal 't_a_253+slope' peakVal
+ t_a_254 peakVal 't_a_254+slope' baseVal
+ t_a_255 baseVal 't_a_255+slope' peakVal
+ t_a_256 peakVal 't_a_256+slope' baseVal
+ t_a_257 baseVal 't_a_257+slope' peakVal
+ t_a_258 peakVal 't_a_258+slope' baseVal
+ t_a_259 baseVal 't_a_259+slope' peakVal
+ t_a_260 peakVal 't_a_260+slope' baseVal
+ t_a_261 baseVal 't_a_261+slope' peakVal
+ t_a_262 peakVal 't_a_262+slope' baseVal
+ t_a_263 baseVal 't_a_263+slope' peakVal
+ t_a_264 peakVal 't_a_264+slope' baseVal
+ t_a_265 baseVal 't_a_265+slope' peakVal
+ t_a_266 peakVal 't_a_266+slope' baseVal
+ t_a_267 baseVal 't_a_267+slope' peakVal
+ t_a_268 peakVal 't_a_268+slope' baseVal
+ t_a_269 baseVal 't_a_269+slope' peakVal
+ t_a_270 peakVal 't_a_270+slope' baseVal
+ t_a_271 baseVal 't_a_271+slope' peakVal
+ t_a_272 peakVal 't_a_272+slope' baseVal
+ t_a_273 baseVal 't_a_273+slope' peakVal
+ t_a_274 peakVal 't_a_274+slope' baseVal
+ t_a_275 baseVal 't_a_275+slope' peakVal
+ t_a_276 peakVal 't_a_276+slope' baseVal
+ t_a_277 baseVal 't_a_277+slope' peakVal
+ t_a_278 peakVal 't_a_278+slope' baseVal
+ t_a_279 baseVal 't_a_279+slope' peakVal
+ t_a_280 peakVal 't_a_280+slope' baseVal
+ t_a_281 baseVal 't_a_281+slope' peakVal
+ t_a_282 peakVal 't_a_282+slope' baseVal
+ t_a_283 baseVal 't_a_283+slope' peakVal
+ t_a_284 peakVal 't_a_284+slope' baseVal
+ t_a_285 baseVal 't_a_285+slope' peakVal
+ t_a_286 peakVal 't_a_286+slope' baseVal
+ t_a_287 baseVal 't_a_287+slope' peakVal
+ t_a_288 peakVal 't_a_288+slope' baseVal
+ t_a_289 baseVal 't_a_289+slope' peakVal
+ t_a_290 peakVal 't_a_290+slope' baseVal
+ t_a_291 baseVal 't_a_291+slope' peakVal
+ t_a_292 peakVal 't_a_292+slope' baseVal
+ t_a_293 baseVal 't_a_293+slope' peakVal
+ t_a_294 peakVal 't_a_294+slope' baseVal
+ t_a_295 baseVal 't_a_295+slope' peakVal
+ t_a_296 peakVal 't_a_296+slope' baseVal
+ t_a_297 baseVal 't_a_297+slope' peakVal
+ t_a_298 peakVal 't_a_298+slope' baseVal
+ t_a_299 baseVal 't_a_299+slope' peakVal
+ t_a_300 peakVal 't_a_300+slope' baseVal
+ t_a_301 baseVal 't_a_301+slope' peakVal
+ t_a_302 peakVal 't_a_302+slope' baseVal
+ t_a_303 baseVal 't_a_303+slope' peakVal
+ t_a_304 peakVal 't_a_304+slope' baseVal
+ t_a_305 baseVal 't_a_305+slope' peakVal
+ t_a_306 peakVal 't_a_306+slope' baseVal
+ t_a_307 baseVal 't_a_307+slope' peakVal
+ t_a_308 peakVal 't_a_308+slope' baseVal
+ t_a_309 baseVal 't_a_309+slope' peakVal
+ t_a_310 peakVal 't_a_310+slope' baseVal
+ t_a_311 baseVal 't_a_311+slope' peakVal
+ t_a_312 peakVal 't_a_312+slope' baseVal
+ t_a_313 baseVal 't_a_313+slope' peakVal
+ t_a_314 peakVal 't_a_314+slope' baseVal
+ t_a_315 baseVal 't_a_315+slope' peakVal
+ t_a_316 peakVal 't_a_316+slope' baseVal
+ t_a_317 baseVal 't_a_317+slope' peakVal
+ t_a_318 peakVal 't_a_318+slope' baseVal
+ t_a_319 baseVal 't_a_319+slope' peakVal
+ t_a_320 peakVal 't_a_320+slope' baseVal
+ t_a_321 baseVal 't_a_321+slope' peakVal
+ t_a_322 peakVal 't_a_322+slope' baseVal
+ t_a_323 baseVal 't_a_323+slope' peakVal
+ t_a_324 peakVal 't_a_324+slope' baseVal
+ t_a_325 baseVal 't_a_325+slope' peakVal
+ t_a_326 peakVal 't_a_326+slope' baseVal
+ t_a_327 baseVal 't_a_327+slope' peakVal
+ t_a_328 peakVal 't_a_328+slope' baseVal
+ t_a_329 baseVal 't_a_329+slope' peakVal
+ t_a_330 peakVal 't_a_330+slope' baseVal
+ t_a_331 baseVal 't_a_331+slope' peakVal
+ t_a_332 peakVal 't_a_332+slope' baseVal
+ t_a_333 baseVal 't_a_333+slope' peakVal
+ t_a_334 peakVal 't_a_334+slope' baseVal
+ t_a_335 baseVal 't_a_335+slope' peakVal
+ t_a_336 peakVal 't_a_336+slope' baseVal
+ t_a_337 baseVal 't_a_337+slope' peakVal
+ t_a_338 peakVal 't_a_338+slope' baseVal
+ t_a_339 baseVal 't_a_339+slope' peakVal
+ t_a_340 peakVal 't_a_340+slope' baseVal
+ t_a_341 baseVal 't_a_341+slope' peakVal
+ t_a_342 peakVal 't_a_342+slope' baseVal
+ t_a_343 baseVal 't_a_343+slope' peakVal
+ t_a_344 peakVal 't_a_344+slope' baseVal
+ t_a_345 baseVal 't_a_345+slope' peakVal
+ t_a_346 peakVal 't_a_346+slope' baseVal
+ t_a_347 baseVal 't_a_347+slope' peakVal
+ t_a_348 peakVal 't_a_348+slope' baseVal
+ t_a_349 baseVal 't_a_349+slope' peakVal
+ t_a_350 peakVal 't_a_350+slope' baseVal
+ t_a_351 baseVal 't_a_351+slope' peakVal
+ t_a_352 peakVal 't_a_352+slope' baseVal
+ t_a_353 baseVal 't_a_353+slope' peakVal
+ t_a_354 peakVal 't_a_354+slope' baseVal
+ t_a_355 baseVal 't_a_355+slope' peakVal
+ t_a_356 peakVal 't_a_356+slope' baseVal
+ t_a_357 baseVal 't_a_357+slope' peakVal
+ t_a_358 peakVal 't_a_358+slope' baseVal
+ t_a_359 baseVal 't_a_359+slope' peakVal
+ t_a_360 peakVal 't_a_360+slope' baseVal
+ t_a_361 baseVal 't_a_361+slope' peakVal
+ t_a_362 peakVal 't_a_362+slope' baseVal
+ t_a_363 baseVal 't_a_363+slope' peakVal
+ t_a_364 peakVal 't_a_364+slope' baseVal
+ t_a_365 baseVal 't_a_365+slope' peakVal
+ t_a_366 peakVal 't_a_366+slope' baseVal
+ t_a_367 baseVal 't_a_367+slope' peakVal
+ t_a_368 peakVal 't_a_368+slope' baseVal
+ t_a_369 baseVal 't_a_369+slope' peakVal
+ t_a_370 peakVal 't_a_370+slope' baseVal
+ t_a_371 baseVal 't_a_371+slope' peakVal
+ t_a_372 peakVal 't_a_372+slope' baseVal
+ t_a_373 baseVal 't_a_373+slope' peakVal
+ t_a_374 peakVal 't_a_374+slope' baseVal
+ t_a_375 baseVal 't_a_375+slope' peakVal
+ t_a_376 peakVal 't_a_376+slope' baseVal
+ t_a_377 baseVal 't_a_377+slope' peakVal
+ t_a_378 peakVal 't_a_378+slope' baseVal
+ t_a_379 baseVal 't_a_379+slope' peakVal
+ t_a_380 peakVal 't_a_380+slope' baseVal
+ t_a_381 baseVal 't_a_381+slope' peakVal
+ t_a_382 peakVal 't_a_382+slope' baseVal
+ t_a_383 baseVal 't_a_383+slope' peakVal
+ t_a_384 peakVal 't_a_384+slope' baseVal
+ t_a_385 baseVal 't_a_385+slope' peakVal
+ t_a_386 peakVal 't_a_386+slope' baseVal
+ t_a_387 baseVal 't_a_387+slope' peakVal
+ t_a_388 peakVal 't_a_388+slope' baseVal
+ t_a_389 baseVal 't_a_389+slope' peakVal
+ t_a_390 peakVal 't_a_390+slope' baseVal
+ t_a_391 baseVal 't_a_391+slope' peakVal
+ t_a_392 peakVal 't_a_392+slope' baseVal
+ t_a_393 baseVal 't_a_393+slope' peakVal
+ t_a_394 peakVal 't_a_394+slope' baseVal
+ t_a_395 baseVal 't_a_395+slope' peakVal
+ t_a_396 peakVal 't_a_396+slope' baseVal
+ t_a_397 baseVal 't_a_397+slope' peakVal
+ t_a_398 peakVal 't_a_398+slope' baseVal
+ t_a_399 baseVal 't_a_399+slope' peakVal
+ t_a_400 peakVal 't_a_400+slope' baseVal
+ t_a_401 baseVal 't_a_401+slope' peakVal
+ t_a_402 peakVal 't_a_402+slope' baseVal
+ t_a_403 baseVal 't_a_403+slope' peakVal
+ t_a_404 peakVal 't_a_404+slope' baseVal
+ t_a_405 baseVal 't_a_405+slope' peakVal
+ t_a_406 peakVal 't_a_406+slope' baseVal
+ t_a_407 baseVal 't_a_407+slope' peakVal
+ t_a_408 peakVal 't_a_408+slope' baseVal
+ t_a_409 baseVal 't_a_409+slope' peakVal
+ t_a_410 peakVal 't_a_410+slope' baseVal
+ t_a_411 baseVal 't_a_411+slope' peakVal
+ t_a_412 peakVal 't_a_412+slope' baseVal
+ t_a_413 baseVal 't_a_413+slope' peakVal
+ t_a_414 peakVal 't_a_414+slope' baseVal
+ t_a_415 baseVal 't_a_415+slope' peakVal
+ t_a_416 peakVal 't_a_416+slope' baseVal
+ t_a_417 baseVal 't_a_417+slope' peakVal
+ t_a_418 peakVal 't_a_418+slope' baseVal
+ t_a_419 baseVal 't_a_419+slope' peakVal
+ t_a_420 peakVal 't_a_420+slope' baseVal
+ t_a_421 baseVal 't_a_421+slope' peakVal
+ t_a_422 peakVal 't_a_422+slope' baseVal
+ t_a_423 baseVal 't_a_423+slope' peakVal
+ t_a_424 peakVal 't_a_424+slope' baseVal
+ t_a_425 baseVal 't_a_425+slope' peakVal
+ t_a_426 peakVal 't_a_426+slope' baseVal
+ t_a_427 baseVal 't_a_427+slope' peakVal
+ t_a_428 peakVal 't_a_428+slope' baseVal
+ t_a_429 baseVal 't_a_429+slope' peakVal
+ t_a_430 peakVal 't_a_430+slope' baseVal
+ t_a_431 baseVal 't_a_431+slope' peakVal
+ t_a_432 peakVal 't_a_432+slope' baseVal
+ t_a_433 baseVal 't_a_433+slope' peakVal
+ t_a_434 peakVal 't_a_434+slope' baseVal
+ t_a_435 baseVal 't_a_435+slope' peakVal
+ t_a_436 peakVal 't_a_436+slope' baseVal
+ t_a_437 baseVal 't_a_437+slope' peakVal
+ t_a_438 peakVal 't_a_438+slope' baseVal
+ t_a_439 baseVal 't_a_439+slope' peakVal
+ t_a_440 peakVal 't_a_440+slope' baseVal
+ t_a_441 baseVal 't_a_441+slope' peakVal
+ t_a_442 peakVal 't_a_442+slope' baseVal
+ t_a_443 baseVal 't_a_443+slope' peakVal
+ t_a_444 peakVal 't_a_444+slope' baseVal
+ t_a_445 baseVal 't_a_445+slope' peakVal
+ t_a_446 peakVal 't_a_446+slope' baseVal
+ t_a_447 baseVal 't_a_447+slope' peakVal
+ t_a_448 peakVal 't_a_448+slope' baseVal
+ t_a_449 baseVal 't_a_449+slope' peakVal
+ t_a_450 peakVal 't_a_450+slope' baseVal
+ t_a_451 baseVal 't_a_451+slope' peakVal
+ t_a_452 peakVal 't_a_452+slope' baseVal
+ t_a_453 baseVal 't_a_453+slope' peakVal
+ t_a_454 peakVal 't_a_454+slope' baseVal
+ t_a_455 baseVal 't_a_455+slope' peakVal
+ t_a_456 peakVal 't_a_456+slope' baseVal
+ t_a_457 baseVal 't_a_457+slope' peakVal
+ t_a_458 peakVal 't_a_458+slope' baseVal
+ t_a_459 baseVal 't_a_459+slope' peakVal
+ t_a_460 peakVal 't_a_460+slope' baseVal
+ t_a_461 baseVal 't_a_461+slope' peakVal
+ t_a_462 peakVal 't_a_462+slope' baseVal
+ t_a_463 baseVal 't_a_463+slope' peakVal
+ t_a_464 peakVal 't_a_464+slope' baseVal
+ t_a_465 baseVal 't_a_465+slope' peakVal
+ t_a_466 peakVal 't_a_466+slope' baseVal
+ t_a_467 baseVal 't_a_467+slope' peakVal
+ t_a_468 peakVal 't_a_468+slope' baseVal
+ t_a_469 baseVal 't_a_469+slope' peakVal
+ t_a_470 peakVal 't_a_470+slope' baseVal
+ t_a_471 baseVal 't_a_471+slope' peakVal
+ t_a_472 peakVal 't_a_472+slope' baseVal
+ t_a_473 baseVal 't_a_473+slope' peakVal
+ t_a_474 peakVal 't_a_474+slope' baseVal
+ t_a_475 baseVal 't_a_475+slope' peakVal
+ t_a_476 peakVal 't_a_476+slope' baseVal
+ t_a_477 baseVal 't_a_477+slope' peakVal
+ t_a_478 peakVal 't_a_478+slope' baseVal
+ t_a_479 baseVal 't_a_479+slope' peakVal
+ t_a_480 peakVal 't_a_480+slope' baseVal
+ t_a_481 baseVal 't_a_481+slope' peakVal
+ t_a_482 peakVal 't_a_482+slope' baseVal
+ t_a_483 baseVal 't_a_483+slope' peakVal
+ t_a_484 peakVal 't_a_484+slope' baseVal
+ t_a_485 baseVal 't_a_485+slope' peakVal
+ t_a_486 peakVal 't_a_486+slope' baseVal
+ t_a_487 baseVal 't_a_487+slope' peakVal
+ t_a_488 peakVal 't_a_488+slope' baseVal
+ t_a_489 baseVal 't_a_489+slope' peakVal
+ t_a_490 peakVal 't_a_490+slope' baseVal
+ t_a_491 baseVal 't_a_491+slope' peakVal
+ t_a_492 peakVal 't_a_492+slope' baseVal
+ t_a_493 baseVal 't_a_493+slope' peakVal
+ t_a_494 peakVal 't_a_494+slope' baseVal
+ t_a_495 baseVal 't_a_495+slope' peakVal
+ t_a_496 peakVal 't_a_496+slope' baseVal
+ t_a_497 baseVal 't_a_497+slope' peakVal
+ t_a_498 peakVal 't_a_498+slope' baseVal
+ t_a_499 baseVal 't_a_499+slope' peakVal
+ t_a_500 peakVal 't_a_500+slope' baseVal
+ t_a_501 baseVal 't_a_501+slope' peakVal
+ t_a_502 peakVal 't_a_502+slope' baseVal
+ t_a_503 baseVal 't_a_503+slope' peakVal
+ t_a_504 peakVal 't_a_504+slope' baseVal
+ t_a_505 baseVal 't_a_505+slope' peakVal
+ t_a_506 peakVal 't_a_506+slope' baseVal
+ t_a_507 baseVal 't_a_507+slope' peakVal
+ t_a_508 peakVal 't_a_508+slope' baseVal
+ t_a_509 baseVal 't_a_509+slope' peakVal
+ t_a_510 peakVal 't_a_510+slope' baseVal
+ t_a_511 baseVal 't_a_511+slope' peakVal
+ t_a_512 peakVal 't_a_512+slope' baseVal
+ t_a_513 baseVal 't_a_513+slope' peakVal
+ t_a_514 peakVal 't_a_514+slope' baseVal
+ t_a_515 baseVal 't_a_515+slope' peakVal
+ t_a_516 peakVal 't_a_516+slope' baseVal
+ t_a_517 baseVal 't_a_517+slope' peakVal
+ t_a_518 peakVal 't_a_518+slope' baseVal
+ t_a_519 baseVal 't_a_519+slope' peakVal
+ t_a_520 peakVal 't_a_520+slope' baseVal
+ t_a_521 baseVal 't_a_521+slope' peakVal
+ t_a_522 peakVal 't_a_522+slope' baseVal
+ t_a_523 baseVal 't_a_523+slope' peakVal
+ t_a_524 peakVal 't_a_524+slope' baseVal
+ t_a_525 baseVal 't_a_525+slope' peakVal
+ t_a_526 peakVal 't_a_526+slope' baseVal
+ t_a_527 baseVal 't_a_527+slope' peakVal
+ t_a_528 peakVal 't_a_528+slope' baseVal
+ t_a_529 baseVal 't_a_529+slope' peakVal
+ t_a_530 peakVal 't_a_530+slope' baseVal
+ t_a_531 baseVal 't_a_531+slope' peakVal
+ t_a_532 peakVal 't_a_532+slope' baseVal
+ t_a_533 baseVal 't_a_533+slope' peakVal
+ t_a_534 peakVal 't_a_534+slope' baseVal
+ t_a_535 baseVal 't_a_535+slope' peakVal
+ t_a_536 peakVal 't_a_536+slope' baseVal
+ t_a_537 baseVal 't_a_537+slope' peakVal
+ t_a_538 peakVal 't_a_538+slope' baseVal
+ t_a_539 baseVal 't_a_539+slope' peakVal
+ t_a_540 peakVal 't_a_540+slope' baseVal
+ t_a_541 baseVal 't_a_541+slope' peakVal
+ t_a_542 peakVal 't_a_542+slope' baseVal
+ t_a_543 baseVal 't_a_543+slope' peakVal
+ t_a_544 peakVal 't_a_544+slope' baseVal
+ t_a_545 baseVal 't_a_545+slope' peakVal
+ t_a_546 peakVal 't_a_546+slope' baseVal
+ t_a_547 baseVal 't_a_547+slope' peakVal
+ t_a_548 peakVal 't_a_548+slope' baseVal
+ t_a_549 baseVal 't_a_549+slope' peakVal
+ t_a_550 peakVal 't_a_550+slope' baseVal
+ t_a_551 baseVal 't_a_551+slope' peakVal
+ t_a_552 peakVal 't_a_552+slope' baseVal
+ t_a_553 baseVal 't_a_553+slope' peakVal
+ t_a_554 peakVal 't_a_554+slope' baseVal
+ t_a_555 baseVal 't_a_555+slope' peakVal
+ t_a_556 peakVal 't_a_556+slope' baseVal
+ t_a_557 baseVal 't_a_557+slope' peakVal
+ t_a_558 peakVal 't_a_558+slope' baseVal
+ t_a_559 baseVal 't_a_559+slope' peakVal
+ t_a_560 peakVal 't_a_560+slope' baseVal
+ t_a_561 baseVal 't_a_561+slope' peakVal
+ t_a_562 peakVal 't_a_562+slope' baseVal
+ t_a_563 baseVal 't_a_563+slope' peakVal
+ t_a_564 peakVal 't_a_564+slope' baseVal
+ t_a_565 baseVal 't_a_565+slope' peakVal
+ t_a_566 peakVal 't_a_566+slope' baseVal
+ t_a_567 baseVal 't_a_567+slope' peakVal
+ t_a_568 peakVal 't_a_568+slope' baseVal
+ t_a_569 baseVal 't_a_569+slope' peakVal
+ t_a_570 peakVal 't_a_570+slope' baseVal
+ t_a_571 baseVal 't_a_571+slope' peakVal
+ t_a_572 peakVal 't_a_572+slope' baseVal
+ t_a_573 baseVal 't_a_573+slope' peakVal
+ t_a_574 peakVal 't_a_574+slope' baseVal
+ t_a_575 baseVal 't_a_575+slope' peakVal
+ t_a_576 peakVal 't_a_576+slope' baseVal
+ t_a_577 baseVal 't_a_577+slope' peakVal
+ t_a_578 peakVal 't_a_578+slope' baseVal
+ t_a_579 baseVal 't_a_579+slope' peakVal
+ t_a_580 peakVal 't_a_580+slope' baseVal
+ t_a_581 baseVal 't_a_581+slope' peakVal
+ t_a_582 peakVal 't_a_582+slope' baseVal
+ t_a_583 baseVal 't_a_583+slope' peakVal
+ t_a_584 peakVal 't_a_584+slope' baseVal
+ t_a_585 baseVal 't_a_585+slope' peakVal
+ t_a_586 peakVal 't_a_586+slope' baseVal
+ t_a_587 baseVal 't_a_587+slope' peakVal
+ t_a_588 peakVal 't_a_588+slope' baseVal
+ t_a_589 baseVal 't_a_589+slope' peakVal
+ t_a_590 peakVal 't_a_590+slope' baseVal
+ t_a_591 baseVal 't_a_591+slope' peakVal
+ t_a_592 peakVal 't_a_592+slope' baseVal
+ t_a_593 baseVal 't_a_593+slope' peakVal
+ t_a_594 peakVal 't_a_594+slope' baseVal
+ t_a_595 baseVal 't_a_595+slope' peakVal
+ t_a_596 peakVal 't_a_596+slope' baseVal
+ t_a_597 baseVal 't_a_597+slope' peakVal
+ t_a_598 peakVal 't_a_598+slope' baseVal
+ t_a_599 baseVal 't_a_599+slope' peakVal
+ t_a_600 peakVal 't_a_600+slope' baseVal
+ t_a_601 baseVal 't_a_601+slope' peakVal
+ t_a_602 peakVal 't_a_602+slope' baseVal
+ t_a_603 baseVal 't_a_603+slope' peakVal
+ t_a_604 peakVal 't_a_604+slope' baseVal
+ t_a_605 baseVal 't_a_605+slope' peakVal
+ t_a_606 peakVal 't_a_606+slope' baseVal
+ t_a_607 baseVal 't_a_607+slope' peakVal
+ t_a_608 peakVal 't_a_608+slope' baseVal
+ t_a_609 baseVal 't_a_609+slope' peakVal
+ t_a_610 peakVal 't_a_610+slope' baseVal
+ t_a_611 baseVal 't_a_611+slope' peakVal
+ t_a_612 peakVal 't_a_612+slope' baseVal
+ t_a_613 baseVal 't_a_613+slope' peakVal
+ t_a_614 peakVal 't_a_614+slope' baseVal
+ t_a_615 baseVal 't_a_615+slope' peakVal
+ t_a_616 peakVal 't_a_616+slope' baseVal
+ t_a_617 baseVal 't_a_617+slope' peakVal
+ t_a_618 peakVal 't_a_618+slope' baseVal
+ t_a_619 baseVal 't_a_619+slope' peakVal
+ t_a_620 peakVal 't_a_620+slope' baseVal
+ t_a_621 baseVal 't_a_621+slope' peakVal
+ t_a_622 peakVal 't_a_622+slope' baseVal
+ t_a_623 baseVal 't_a_623+slope' peakVal
+ t_a_624 peakVal 't_a_624+slope' baseVal
+ t_a_625 baseVal 't_a_625+slope' peakVal
+ t_a_626 peakVal 't_a_626+slope' baseVal
+ t_a_627 baseVal 't_a_627+slope' peakVal
+ t_a_628 peakVal 't_a_628+slope' baseVal
+ t_a_629 baseVal 't_a_629+slope' peakVal
+ t_a_630 peakVal 't_a_630+slope' baseVal
+ t_a_631 baseVal 't_a_631+slope' peakVal
+ t_a_632 peakVal 't_a_632+slope' baseVal
+ t_a_633 baseVal 't_a_633+slope' peakVal
+ t_a_634 peakVal 't_a_634+slope' baseVal
+ t_a_635 baseVal 't_a_635+slope' peakVal
+ t_a_636 peakVal 't_a_636+slope' baseVal
+ t_a_637 baseVal 't_a_637+slope' peakVal
+ t_a_638 peakVal 't_a_638+slope' baseVal
+ t_a_639 baseVal 't_a_639+slope' peakVal
+ t_a_640 peakVal 't_a_640+slope' baseVal
+ t_a_641 baseVal 't_a_641+slope' peakVal
+ t_a_642 peakVal 't_a_642+slope' baseVal
+ t_a_643 baseVal 't_a_643+slope' peakVal
+ t_a_644 peakVal 't_a_644+slope' baseVal
+ t_a_645 baseVal 't_a_645+slope' peakVal
+ t_a_646 peakVal 't_a_646+slope' baseVal
+ t_a_647 baseVal 't_a_647+slope' peakVal
+ t_a_648 peakVal 't_a_648+slope' baseVal
+ t_a_649 baseVal 't_a_649+slope' peakVal
+ t_a_650 peakVal 't_a_650+slope' baseVal
+ t_a_651 baseVal 't_a_651+slope' peakVal
+ t_a_652 peakVal 't_a_652+slope' baseVal
+ t_a_653 baseVal 't_a_653+slope' peakVal
+ t_a_654 peakVal 't_a_654+slope' baseVal
+ t_a_655 baseVal 't_a_655+slope' peakVal
+ t_a_656 peakVal 't_a_656+slope' baseVal
+ t_a_657 baseVal 't_a_657+slope' peakVal
+ t_a_658 peakVal 't_a_658+slope' baseVal
+ t_a_659 baseVal 't_a_659+slope' peakVal
+ t_a_660 peakVal 't_a_660+slope' baseVal
+ t_a_661 baseVal 't_a_661+slope' peakVal
+ t_a_662 peakVal 't_a_662+slope' baseVal
+ t_a_663 baseVal 't_a_663+slope' peakVal
+ t_a_664 peakVal 't_a_664+slope' baseVal
+ t_a_665 baseVal 't_a_665+slope' peakVal
+ t_a_666 peakVal 't_a_666+slope' baseVal
+ t_a_667 baseVal 't_a_667+slope' peakVal
+ t_a_668 peakVal 't_a_668+slope' baseVal
+ t_a_669 baseVal 't_a_669+slope' peakVal
+ t_a_670 peakVal 't_a_670+slope' baseVal
+ t_a_671 baseVal 't_a_671+slope' peakVal
+ t_a_672 peakVal 't_a_672+slope' baseVal
+ t_a_673 baseVal 't_a_673+slope' peakVal
+ t_a_674 peakVal 't_a_674+slope' baseVal
+ t_a_675 baseVal 't_a_675+slope' peakVal
+ t_a_676 peakVal 't_a_676+slope' baseVal
+ t_a_677 baseVal 't_a_677+slope' peakVal
+ t_a_678 peakVal 't_a_678+slope' baseVal
+ t_a_679 baseVal 't_a_679+slope' peakVal
+ t_a_680 peakVal 't_a_680+slope' baseVal
+ t_a_681 baseVal 't_a_681+slope' peakVal
+ t_a_682 peakVal 't_a_682+slope' baseVal
+ t_a_683 baseVal 't_a_683+slope' peakVal
+ t_a_684 peakVal 't_a_684+slope' baseVal
+ t_a_685 baseVal 't_a_685+slope' peakVal
+ t_a_686 peakVal 't_a_686+slope' baseVal
+ t_a_687 baseVal 't_a_687+slope' peakVal
+ t_a_688 peakVal 't_a_688+slope' baseVal
+ t_a_689 baseVal 't_a_689+slope' peakVal
+ t_a_690 peakVal 't_a_690+slope' baseVal
+ t_a_691 baseVal 't_a_691+slope' peakVal
+ t_a_692 peakVal 't_a_692+slope' baseVal
+ t_a_693 baseVal 't_a_693+slope' peakVal
+ t_a_694 peakVal 't_a_694+slope' baseVal
+ t_a_695 baseVal 't_a_695+slope' peakVal
+ t_a_696 peakVal 't_a_696+slope' baseVal
+ t_a_697 baseVal 't_a_697+slope' peakVal
+ t_a_698 peakVal 't_a_698+slope' baseVal
+ t_a_699 baseVal 't_a_699+slope' peakVal
+ t_a_700 peakVal 't_a_700+slope' baseVal
+ t_a_701 baseVal 't_a_701+slope' peakVal
+ t_a_702 peakVal 't_a_702+slope' baseVal
+ t_a_703 baseVal 't_a_703+slope' peakVal
+ t_a_704 peakVal 't_a_704+slope' baseVal
+ t_a_705 baseVal 't_a_705+slope' peakVal
+ t_a_706 peakVal 't_a_706+slope' baseVal
+ t_a_707 baseVal 't_a_707+slope' peakVal
+ t_a_708 peakVal 't_a_708+slope' baseVal
+ t_a_709 baseVal 't_a_709+slope' peakVal
+ t_a_710 peakVal 't_a_710+slope' baseVal
+ t_a_711 baseVal 't_a_711+slope' peakVal
+ t_a_712 peakVal 't_a_712+slope' baseVal
+ t_a_713 baseVal 't_a_713+slope' peakVal
+ t_a_714 peakVal 't_a_714+slope' baseVal
+ t_a_715 baseVal 't_a_715+slope' peakVal
+ t_a_716 peakVal 't_a_716+slope' baseVal
+ t_a_717 baseVal 't_a_717+slope' peakVal
+ t_a_718 peakVal 't_a_718+slope' baseVal
+ t_a_719 baseVal 't_a_719+slope' peakVal
+ t_a_720 peakVal 't_a_720+slope' baseVal
+ t_a_721 baseVal 't_a_721+slope' peakVal
+ t_a_722 peakVal 't_a_722+slope' baseVal
+ t_a_723 baseVal 't_a_723+slope' peakVal
+ t_a_724 peakVal 't_a_724+slope' baseVal
+ t_a_725 baseVal 't_a_725+slope' peakVal
+ t_a_726 peakVal 't_a_726+slope' baseVal
+ t_a_727 baseVal 't_a_727+slope' peakVal
+ t_a_728 peakVal 't_a_728+slope' baseVal
+ t_a_729 baseVal 't_a_729+slope' peakVal
+ t_a_730 peakVal 't_a_730+slope' baseVal
+ t_a_731 baseVal 't_a_731+slope' peakVal
+ t_a_732 peakVal 't_a_732+slope' baseVal
+ t_a_733 baseVal 't_a_733+slope' peakVal
+ t_a_734 peakVal 't_a_734+slope' baseVal
+ t_a_735 baseVal 't_a_735+slope' peakVal
+ t_a_736 peakVal 't_a_736+slope' baseVal
+ t_a_737 baseVal 't_a_737+slope' peakVal
+ t_a_738 peakVal 't_a_738+slope' baseVal
+ t_a_739 baseVal 't_a_739+slope' peakVal
+ t_a_740 peakVal 't_a_740+slope' baseVal
+ t_a_741 baseVal 't_a_741+slope' peakVal
+ t_a_742 peakVal 't_a_742+slope' baseVal
+ t_a_743 baseVal 't_a_743+slope' peakVal
+ t_a_744 peakVal 't_a_744+slope' baseVal
+ t_a_745 baseVal 't_a_745+slope' peakVal
+ t_a_746 peakVal 't_a_746+slope' baseVal
+ t_a_747 baseVal 't_a_747+slope' peakVal
+ t_a_748 peakVal 't_a_748+slope' baseVal
+ t_a_749 baseVal 't_a_749+slope' peakVal
+ t_a_750 peakVal 't_a_750+slope' baseVal
+ t_a_751 baseVal 't_a_751+slope' peakVal
+ t_a_752 peakVal 't_a_752+slope' baseVal
+ t_a_753 baseVal 't_a_753+slope' peakVal
+ t_a_754 peakVal 't_a_754+slope' baseVal
+ t_a_755 baseVal 't_a_755+slope' peakVal
+ t_a_756 peakVal 't_a_756+slope' baseVal
+ t_a_757 baseVal 't_a_757+slope' peakVal
+ t_a_758 peakVal 't_a_758+slope' baseVal
+ t_a_759 baseVal 't_a_759+slope' peakVal
+ t_a_760 peakVal 't_a_760+slope' baseVal
+ t_a_761 baseVal 't_a_761+slope' peakVal
+ t_a_762 peakVal 't_a_762+slope' baseVal
+ t_a_763 baseVal 't_a_763+slope' peakVal
+ t_a_764 peakVal 't_a_764+slope' baseVal
+ t_a_765 baseVal 't_a_765+slope' peakVal
+ t_a_766 peakVal 't_a_766+slope' baseVal
+ t_a_767 baseVal 't_a_767+slope' peakVal
+ t_a_768 peakVal 't_a_768+slope' baseVal
+ t_a_769 baseVal 't_a_769+slope' peakVal
+ t_a_770 peakVal 't_a_770+slope' baseVal
+ t_a_771 baseVal 't_a_771+slope' peakVal
+ t_a_772 peakVal 't_a_772+slope' baseVal
+ t_a_773 baseVal 't_a_773+slope' peakVal
+ t_a_774 peakVal 't_a_774+slope' baseVal
+ t_a_775 baseVal 't_a_775+slope' peakVal
+ t_a_776 peakVal 't_a_776+slope' baseVal
+ t_a_777 baseVal 't_a_777+slope' peakVal
+ t_a_778 peakVal 't_a_778+slope' baseVal
+ t_a_779 baseVal 't_a_779+slope' peakVal
+ t_a_780 peakVal 't_a_780+slope' baseVal
+ t_a_781 baseVal 't_a_781+slope' peakVal
+ t_a_782 peakVal 't_a_782+slope' baseVal
+ t_a_783 baseVal 't_a_783+slope' peakVal
+ t_a_784 peakVal 't_a_784+slope' baseVal
+ t_a_785 baseVal 't_a_785+slope' peakVal
+ t_a_786 peakVal 't_a_786+slope' baseVal
+ t_a_787 baseVal 't_a_787+slope' peakVal
+ t_a_788 peakVal 't_a_788+slope' baseVal
+ t_a_789 baseVal 't_a_789+slope' peakVal
+ t_a_790 peakVal 't_a_790+slope' baseVal
+ t_a_791 baseVal 't_a_791+slope' peakVal
+ t_a_792 peakVal 't_a_792+slope' baseVal
+ t_a_793 baseVal 't_a_793+slope' peakVal
+ t_a_794 peakVal 't_a_794+slope' baseVal
+ t_a_795 baseVal 't_a_795+slope' peakVal
+ t_a_796 peakVal 't_a_796+slope' baseVal
+ t_a_797 baseVal 't_a_797+slope' peakVal
+ t_a_798 peakVal 't_a_798+slope' baseVal
+ t_a_799 baseVal 't_a_799+slope' peakVal



VINB Input_B GND PWL 0ns baseVal t_init0 baseVal 't_init0+slope' peakVal t_init1 peakVal 't_init1+slope' baseVal
+ t_b_0 peakVal 't_b_0+slope' baseVal
+ t_b_1 baseVal 't_b_1+slope' peakVal
+ t_b_2 peakVal 't_b_2+slope' baseVal
+ t_b_3 baseVal 't_b_3+slope' peakVal
+ t_b_4 peakVal 't_b_4+slope' baseVal
+ t_b_5 baseVal 't_b_5+slope' peakVal
+ t_b_6 peakVal 't_b_6+slope' baseVal
+ t_b_7 baseVal 't_b_7+slope' peakVal
+ t_b_8 peakVal 't_b_8+slope' baseVal
+ t_b_9 baseVal 't_b_9+slope' peakVal
+ t_b_10 peakVal 't_b_10+slope' baseVal
+ t_b_11 baseVal 't_b_11+slope' peakVal
+ t_b_12 peakVal 't_b_12+slope' baseVal
+ t_b_13 baseVal 't_b_13+slope' peakVal
+ t_b_14 peakVal 't_b_14+slope' baseVal
+ t_b_15 baseVal 't_b_15+slope' peakVal
+ t_b_16 peakVal 't_b_16+slope' baseVal
+ t_b_17 baseVal 't_b_17+slope' peakVal
+ t_b_18 peakVal 't_b_18+slope' baseVal
+ t_b_19 baseVal 't_b_19+slope' peakVal
+ t_b_20 peakVal 't_b_20+slope' baseVal
+ t_b_21 baseVal 't_b_21+slope' peakVal
+ t_b_22 peakVal 't_b_22+slope' baseVal
+ t_b_23 baseVal 't_b_23+slope' peakVal
+ t_b_24 peakVal 't_b_24+slope' baseVal
+ t_b_25 baseVal 't_b_25+slope' peakVal
+ t_b_26 peakVal 't_b_26+slope' baseVal
+ t_b_27 baseVal 't_b_27+slope' peakVal
+ t_b_28 peakVal 't_b_28+slope' baseVal
+ t_b_29 baseVal 't_b_29+slope' peakVal
+ t_b_30 peakVal 't_b_30+slope' baseVal
+ t_b_31 baseVal 't_b_31+slope' peakVal
+ t_b_32 peakVal 't_b_32+slope' baseVal
+ t_b_33 baseVal 't_b_33+slope' peakVal
+ t_b_34 peakVal 't_b_34+slope' baseVal
+ t_b_35 baseVal 't_b_35+slope' peakVal
+ t_b_36 peakVal 't_b_36+slope' baseVal
+ t_b_37 baseVal 't_b_37+slope' peakVal
+ t_b_38 peakVal 't_b_38+slope' baseVal
+ t_b_39 baseVal 't_b_39+slope' peakVal
+ t_b_40 peakVal 't_b_40+slope' baseVal
+ t_b_41 baseVal 't_b_41+slope' peakVal
+ t_b_42 peakVal 't_b_42+slope' baseVal
+ t_b_43 baseVal 't_b_43+slope' peakVal
+ t_b_44 peakVal 't_b_44+slope' baseVal
+ t_b_45 baseVal 't_b_45+slope' peakVal
+ t_b_46 peakVal 't_b_46+slope' baseVal
+ t_b_47 baseVal 't_b_47+slope' peakVal
+ t_b_48 peakVal 't_b_48+slope' baseVal
+ t_b_49 baseVal 't_b_49+slope' peakVal
+ t_b_50 peakVal 't_b_50+slope' baseVal
+ t_b_51 baseVal 't_b_51+slope' peakVal
+ t_b_52 peakVal 't_b_52+slope' baseVal
+ t_b_53 baseVal 't_b_53+slope' peakVal
+ t_b_54 peakVal 't_b_54+slope' baseVal
+ t_b_55 baseVal 't_b_55+slope' peakVal
+ t_b_56 peakVal 't_b_56+slope' baseVal
+ t_b_57 baseVal 't_b_57+slope' peakVal
+ t_b_58 peakVal 't_b_58+slope' baseVal
+ t_b_59 baseVal 't_b_59+slope' peakVal
+ t_b_60 peakVal 't_b_60+slope' baseVal
+ t_b_61 baseVal 't_b_61+slope' peakVal
+ t_b_62 peakVal 't_b_62+slope' baseVal
+ t_b_63 baseVal 't_b_63+slope' peakVal
+ t_b_64 peakVal 't_b_64+slope' baseVal
+ t_b_65 baseVal 't_b_65+slope' peakVal
+ t_b_66 peakVal 't_b_66+slope' baseVal
+ t_b_67 baseVal 't_b_67+slope' peakVal
+ t_b_68 peakVal 't_b_68+slope' baseVal
+ t_b_69 baseVal 't_b_69+slope' peakVal
+ t_b_70 peakVal 't_b_70+slope' baseVal
+ t_b_71 baseVal 't_b_71+slope' peakVal
+ t_b_72 peakVal 't_b_72+slope' baseVal
+ t_b_73 baseVal 't_b_73+slope' peakVal
+ t_b_74 peakVal 't_b_74+slope' baseVal
+ t_b_75 baseVal 't_b_75+slope' peakVal
+ t_b_76 peakVal 't_b_76+slope' baseVal
+ t_b_77 baseVal 't_b_77+slope' peakVal
+ t_b_78 peakVal 't_b_78+slope' baseVal
+ t_b_79 baseVal 't_b_79+slope' peakVal
+ t_b_80 peakVal 't_b_80+slope' baseVal
+ t_b_81 baseVal 't_b_81+slope' peakVal
+ t_b_82 peakVal 't_b_82+slope' baseVal
+ t_b_83 baseVal 't_b_83+slope' peakVal
+ t_b_84 peakVal 't_b_84+slope' baseVal
+ t_b_85 baseVal 't_b_85+slope' peakVal
+ t_b_86 peakVal 't_b_86+slope' baseVal
+ t_b_87 baseVal 't_b_87+slope' peakVal
+ t_b_88 peakVal 't_b_88+slope' baseVal
+ t_b_89 baseVal 't_b_89+slope' peakVal
+ t_b_90 peakVal 't_b_90+slope' baseVal
+ t_b_91 baseVal 't_b_91+slope' peakVal
+ t_b_92 peakVal 't_b_92+slope' baseVal
+ t_b_93 baseVal 't_b_93+slope' peakVal
+ t_b_94 peakVal 't_b_94+slope' baseVal
+ t_b_95 baseVal 't_b_95+slope' peakVal
+ t_b_96 peakVal 't_b_96+slope' baseVal
+ t_b_97 baseVal 't_b_97+slope' peakVal
+ t_b_98 peakVal 't_b_98+slope' baseVal
+ t_b_99 baseVal 't_b_99+slope' peakVal
+ t_b_100 peakVal 't_b_100+slope' baseVal
+ t_b_101 baseVal 't_b_101+slope' peakVal
+ t_b_102 peakVal 't_b_102+slope' baseVal
+ t_b_103 baseVal 't_b_103+slope' peakVal
+ t_b_104 peakVal 't_b_104+slope' baseVal
+ t_b_105 baseVal 't_b_105+slope' peakVal
+ t_b_106 peakVal 't_b_106+slope' baseVal
+ t_b_107 baseVal 't_b_107+slope' peakVal
+ t_b_108 peakVal 't_b_108+slope' baseVal
+ t_b_109 baseVal 't_b_109+slope' peakVal
+ t_b_110 peakVal 't_b_110+slope' baseVal
+ t_b_111 baseVal 't_b_111+slope' peakVal
+ t_b_112 peakVal 't_b_112+slope' baseVal
+ t_b_113 baseVal 't_b_113+slope' peakVal
+ t_b_114 peakVal 't_b_114+slope' baseVal
+ t_b_115 baseVal 't_b_115+slope' peakVal
+ t_b_116 peakVal 't_b_116+slope' baseVal
+ t_b_117 baseVal 't_b_117+slope' peakVal
+ t_b_118 peakVal 't_b_118+slope' baseVal
+ t_b_119 baseVal 't_b_119+slope' peakVal
+ t_b_120 peakVal 't_b_120+slope' baseVal
+ t_b_121 baseVal 't_b_121+slope' peakVal
+ t_b_122 peakVal 't_b_122+slope' baseVal
+ t_b_123 baseVal 't_b_123+slope' peakVal
+ t_b_124 peakVal 't_b_124+slope' baseVal
+ t_b_125 baseVal 't_b_125+slope' peakVal
+ t_b_126 peakVal 't_b_126+slope' baseVal
+ t_b_127 baseVal 't_b_127+slope' peakVal
+ t_b_128 peakVal 't_b_128+slope' baseVal
+ t_b_129 baseVal 't_b_129+slope' peakVal
+ t_b_130 peakVal 't_b_130+slope' baseVal
+ t_b_131 baseVal 't_b_131+slope' peakVal
+ t_b_132 peakVal 't_b_132+slope' baseVal
+ t_b_133 baseVal 't_b_133+slope' peakVal
+ t_b_134 peakVal 't_b_134+slope' baseVal
+ t_b_135 baseVal 't_b_135+slope' peakVal
+ t_b_136 peakVal 't_b_136+slope' baseVal
+ t_b_137 baseVal 't_b_137+slope' peakVal
+ t_b_138 peakVal 't_b_138+slope' baseVal
+ t_b_139 baseVal 't_b_139+slope' peakVal
+ t_b_140 peakVal 't_b_140+slope' baseVal
+ t_b_141 baseVal 't_b_141+slope' peakVal
+ t_b_142 peakVal 't_b_142+slope' baseVal
+ t_b_143 baseVal 't_b_143+slope' peakVal
+ t_b_144 peakVal 't_b_144+slope' baseVal
+ t_b_145 baseVal 't_b_145+slope' peakVal
+ t_b_146 peakVal 't_b_146+slope' baseVal
+ t_b_147 baseVal 't_b_147+slope' peakVal
+ t_b_148 peakVal 't_b_148+slope' baseVal
+ t_b_149 baseVal 't_b_149+slope' peakVal
+ t_b_150 peakVal 't_b_150+slope' baseVal
+ t_b_151 baseVal 't_b_151+slope' peakVal
+ t_b_152 peakVal 't_b_152+slope' baseVal
+ t_b_153 baseVal 't_b_153+slope' peakVal
+ t_b_154 peakVal 't_b_154+slope' baseVal
+ t_b_155 baseVal 't_b_155+slope' peakVal
+ t_b_156 peakVal 't_b_156+slope' baseVal
+ t_b_157 baseVal 't_b_157+slope' peakVal
+ t_b_158 peakVal 't_b_158+slope' baseVal
+ t_b_159 baseVal 't_b_159+slope' peakVal
+ t_b_160 peakVal 't_b_160+slope' baseVal
+ t_b_161 baseVal 't_b_161+slope' peakVal
+ t_b_162 peakVal 't_b_162+slope' baseVal
+ t_b_163 baseVal 't_b_163+slope' peakVal
+ t_b_164 peakVal 't_b_164+slope' baseVal
+ t_b_165 baseVal 't_b_165+slope' peakVal
+ t_b_166 peakVal 't_b_166+slope' baseVal
+ t_b_167 baseVal 't_b_167+slope' peakVal
+ t_b_168 peakVal 't_b_168+slope' baseVal
+ t_b_169 baseVal 't_b_169+slope' peakVal
+ t_b_170 peakVal 't_b_170+slope' baseVal
+ t_b_171 baseVal 't_b_171+slope' peakVal
+ t_b_172 peakVal 't_b_172+slope' baseVal
+ t_b_173 baseVal 't_b_173+slope' peakVal
+ t_b_174 peakVal 't_b_174+slope' baseVal
+ t_b_175 baseVal 't_b_175+slope' peakVal
+ t_b_176 peakVal 't_b_176+slope' baseVal
+ t_b_177 baseVal 't_b_177+slope' peakVal
+ t_b_178 peakVal 't_b_178+slope' baseVal
+ t_b_179 baseVal 't_b_179+slope' peakVal
+ t_b_180 peakVal 't_b_180+slope' baseVal
+ t_b_181 baseVal 't_b_181+slope' peakVal
+ t_b_182 peakVal 't_b_182+slope' baseVal
+ t_b_183 baseVal 't_b_183+slope' peakVal
+ t_b_184 peakVal 't_b_184+slope' baseVal
+ t_b_185 baseVal 't_b_185+slope' peakVal
+ t_b_186 peakVal 't_b_186+slope' baseVal
+ t_b_187 baseVal 't_b_187+slope' peakVal
+ t_b_188 peakVal 't_b_188+slope' baseVal
+ t_b_189 baseVal 't_b_189+slope' peakVal
+ t_b_190 peakVal 't_b_190+slope' baseVal
+ t_b_191 baseVal 't_b_191+slope' peakVal
+ t_b_192 peakVal 't_b_192+slope' baseVal
+ t_b_193 baseVal 't_b_193+slope' peakVal
+ t_b_194 peakVal 't_b_194+slope' baseVal
+ t_b_195 baseVal 't_b_195+slope' peakVal
+ t_b_196 peakVal 't_b_196+slope' baseVal
+ t_b_197 baseVal 't_b_197+slope' peakVal
+ t_b_198 peakVal 't_b_198+slope' baseVal
+ t_b_199 baseVal 't_b_199+slope' peakVal
+ t_b_200 peakVal 't_b_200+slope' baseVal
+ t_b_201 baseVal 't_b_201+slope' peakVal
+ t_b_202 peakVal 't_b_202+slope' baseVal
+ t_b_203 baseVal 't_b_203+slope' peakVal
+ t_b_204 peakVal 't_b_204+slope' baseVal
+ t_b_205 baseVal 't_b_205+slope' peakVal
+ t_b_206 peakVal 't_b_206+slope' baseVal
+ t_b_207 baseVal 't_b_207+slope' peakVal
+ t_b_208 peakVal 't_b_208+slope' baseVal
+ t_b_209 baseVal 't_b_209+slope' peakVal
+ t_b_210 peakVal 't_b_210+slope' baseVal
+ t_b_211 baseVal 't_b_211+slope' peakVal
+ t_b_212 peakVal 't_b_212+slope' baseVal
+ t_b_213 baseVal 't_b_213+slope' peakVal
+ t_b_214 peakVal 't_b_214+slope' baseVal
+ t_b_215 baseVal 't_b_215+slope' peakVal
+ t_b_216 peakVal 't_b_216+slope' baseVal
+ t_b_217 baseVal 't_b_217+slope' peakVal
+ t_b_218 peakVal 't_b_218+slope' baseVal
+ t_b_219 baseVal 't_b_219+slope' peakVal
+ t_b_220 peakVal 't_b_220+slope' baseVal
+ t_b_221 baseVal 't_b_221+slope' peakVal
+ t_b_222 peakVal 't_b_222+slope' baseVal
+ t_b_223 baseVal 't_b_223+slope' peakVal
+ t_b_224 peakVal 't_b_224+slope' baseVal
+ t_b_225 baseVal 't_b_225+slope' peakVal
+ t_b_226 peakVal 't_b_226+slope' baseVal
+ t_b_227 baseVal 't_b_227+slope' peakVal
+ t_b_228 peakVal 't_b_228+slope' baseVal
+ t_b_229 baseVal 't_b_229+slope' peakVal
+ t_b_230 peakVal 't_b_230+slope' baseVal
+ t_b_231 baseVal 't_b_231+slope' peakVal
+ t_b_232 peakVal 't_b_232+slope' baseVal
+ t_b_233 baseVal 't_b_233+slope' peakVal
+ t_b_234 peakVal 't_b_234+slope' baseVal
+ t_b_235 baseVal 't_b_235+slope' peakVal
+ t_b_236 peakVal 't_b_236+slope' baseVal
+ t_b_237 baseVal 't_b_237+slope' peakVal
+ t_b_238 peakVal 't_b_238+slope' baseVal
+ t_b_239 baseVal 't_b_239+slope' peakVal
+ t_b_240 peakVal 't_b_240+slope' baseVal
+ t_b_241 baseVal 't_b_241+slope' peakVal
+ t_b_242 peakVal 't_b_242+slope' baseVal
+ t_b_243 baseVal 't_b_243+slope' peakVal
+ t_b_244 peakVal 't_b_244+slope' baseVal
+ t_b_245 baseVal 't_b_245+slope' peakVal
+ t_b_246 peakVal 't_b_246+slope' baseVal
+ t_b_247 baseVal 't_b_247+slope' peakVal
+ t_b_248 peakVal 't_b_248+slope' baseVal
+ t_b_249 baseVal 't_b_249+slope' peakVal
+ t_b_250 peakVal 't_b_250+slope' baseVal
+ t_b_251 baseVal 't_b_251+slope' peakVal
+ t_b_252 peakVal 't_b_252+slope' baseVal
+ t_b_253 baseVal 't_b_253+slope' peakVal
+ t_b_254 peakVal 't_b_254+slope' baseVal
+ t_b_255 baseVal 't_b_255+slope' peakVal
+ t_b_256 peakVal 't_b_256+slope' baseVal
+ t_b_257 baseVal 't_b_257+slope' peakVal
+ t_b_258 peakVal 't_b_258+slope' baseVal
+ t_b_259 baseVal 't_b_259+slope' peakVal
+ t_b_260 peakVal 't_b_260+slope' baseVal
+ t_b_261 baseVal 't_b_261+slope' peakVal
+ t_b_262 peakVal 't_b_262+slope' baseVal
+ t_b_263 baseVal 't_b_263+slope' peakVal
+ t_b_264 peakVal 't_b_264+slope' baseVal
+ t_b_265 baseVal 't_b_265+slope' peakVal
+ t_b_266 peakVal 't_b_266+slope' baseVal
+ t_b_267 baseVal 't_b_267+slope' peakVal
+ t_b_268 peakVal 't_b_268+slope' baseVal
+ t_b_269 baseVal 't_b_269+slope' peakVal
+ t_b_270 peakVal 't_b_270+slope' baseVal
+ t_b_271 baseVal 't_b_271+slope' peakVal
+ t_b_272 peakVal 't_b_272+slope' baseVal
+ t_b_273 baseVal 't_b_273+slope' peakVal
+ t_b_274 peakVal 't_b_274+slope' baseVal
+ t_b_275 baseVal 't_b_275+slope' peakVal
+ t_b_276 peakVal 't_b_276+slope' baseVal
+ t_b_277 baseVal 't_b_277+slope' peakVal
+ t_b_278 peakVal 't_b_278+slope' baseVal
+ t_b_279 baseVal 't_b_279+slope' peakVal
+ t_b_280 peakVal 't_b_280+slope' baseVal
+ t_b_281 baseVal 't_b_281+slope' peakVal
+ t_b_282 peakVal 't_b_282+slope' baseVal
+ t_b_283 baseVal 't_b_283+slope' peakVal
+ t_b_284 peakVal 't_b_284+slope' baseVal
+ t_b_285 baseVal 't_b_285+slope' peakVal
+ t_b_286 peakVal 't_b_286+slope' baseVal
+ t_b_287 baseVal 't_b_287+slope' peakVal
+ t_b_288 peakVal 't_b_288+slope' baseVal
+ t_b_289 baseVal 't_b_289+slope' peakVal
+ t_b_290 peakVal 't_b_290+slope' baseVal
+ t_b_291 baseVal 't_b_291+slope' peakVal
+ t_b_292 peakVal 't_b_292+slope' baseVal
+ t_b_293 baseVal 't_b_293+slope' peakVal
+ t_b_294 peakVal 't_b_294+slope' baseVal
+ t_b_295 baseVal 't_b_295+slope' peakVal
+ t_b_296 peakVal 't_b_296+slope' baseVal
+ t_b_297 baseVal 't_b_297+slope' peakVal
+ t_b_298 peakVal 't_b_298+slope' baseVal
+ t_b_299 baseVal 't_b_299+slope' peakVal
+ t_b_300 peakVal 't_b_300+slope' baseVal
+ t_b_301 baseVal 't_b_301+slope' peakVal
+ t_b_302 peakVal 't_b_302+slope' baseVal
+ t_b_303 baseVal 't_b_303+slope' peakVal
+ t_b_304 peakVal 't_b_304+slope' baseVal
+ t_b_305 baseVal 't_b_305+slope' peakVal
+ t_b_306 peakVal 't_b_306+slope' baseVal
+ t_b_307 baseVal 't_b_307+slope' peakVal
+ t_b_308 peakVal 't_b_308+slope' baseVal
+ t_b_309 baseVal 't_b_309+slope' peakVal
+ t_b_310 peakVal 't_b_310+slope' baseVal
+ t_b_311 baseVal 't_b_311+slope' peakVal
+ t_b_312 peakVal 't_b_312+slope' baseVal
+ t_b_313 baseVal 't_b_313+slope' peakVal
+ t_b_314 peakVal 't_b_314+slope' baseVal
+ t_b_315 baseVal 't_b_315+slope' peakVal
+ t_b_316 peakVal 't_b_316+slope' baseVal
+ t_b_317 baseVal 't_b_317+slope' peakVal
+ t_b_318 peakVal 't_b_318+slope' baseVal
+ t_b_319 baseVal 't_b_319+slope' peakVal
+ t_b_320 peakVal 't_b_320+slope' baseVal
+ t_b_321 baseVal 't_b_321+slope' peakVal
+ t_b_322 peakVal 't_b_322+slope' baseVal
+ t_b_323 baseVal 't_b_323+slope' peakVal
+ t_b_324 peakVal 't_b_324+slope' baseVal
+ t_b_325 baseVal 't_b_325+slope' peakVal
+ t_b_326 peakVal 't_b_326+slope' baseVal
+ t_b_327 baseVal 't_b_327+slope' peakVal
+ t_b_328 peakVal 't_b_328+slope' baseVal
+ t_b_329 baseVal 't_b_329+slope' peakVal
+ t_b_330 peakVal 't_b_330+slope' baseVal
+ t_b_331 baseVal 't_b_331+slope' peakVal
+ t_b_332 peakVal 't_b_332+slope' baseVal
+ t_b_333 baseVal 't_b_333+slope' peakVal
+ t_b_334 peakVal 't_b_334+slope' baseVal
+ t_b_335 baseVal 't_b_335+slope' peakVal
+ t_b_336 peakVal 't_b_336+slope' baseVal
+ t_b_337 baseVal 't_b_337+slope' peakVal
+ t_b_338 peakVal 't_b_338+slope' baseVal
+ t_b_339 baseVal 't_b_339+slope' peakVal
+ t_b_340 peakVal 't_b_340+slope' baseVal
+ t_b_341 baseVal 't_b_341+slope' peakVal
+ t_b_342 peakVal 't_b_342+slope' baseVal
+ t_b_343 baseVal 't_b_343+slope' peakVal
+ t_b_344 peakVal 't_b_344+slope' baseVal
+ t_b_345 baseVal 't_b_345+slope' peakVal
+ t_b_346 peakVal 't_b_346+slope' baseVal
+ t_b_347 baseVal 't_b_347+slope' peakVal
+ t_b_348 peakVal 't_b_348+slope' baseVal
+ t_b_349 baseVal 't_b_349+slope' peakVal
+ t_b_350 peakVal 't_b_350+slope' baseVal
+ t_b_351 baseVal 't_b_351+slope' peakVal
+ t_b_352 peakVal 't_b_352+slope' baseVal
+ t_b_353 baseVal 't_b_353+slope' peakVal
+ t_b_354 peakVal 't_b_354+slope' baseVal
+ t_b_355 baseVal 't_b_355+slope' peakVal
+ t_b_356 peakVal 't_b_356+slope' baseVal
+ t_b_357 baseVal 't_b_357+slope' peakVal
+ t_b_358 peakVal 't_b_358+slope' baseVal
+ t_b_359 baseVal 't_b_359+slope' peakVal
+ t_b_360 peakVal 't_b_360+slope' baseVal
+ t_b_361 baseVal 't_b_361+slope' peakVal
+ t_b_362 peakVal 't_b_362+slope' baseVal
+ t_b_363 baseVal 't_b_363+slope' peakVal
+ t_b_364 peakVal 't_b_364+slope' baseVal
+ t_b_365 baseVal 't_b_365+slope' peakVal
+ t_b_366 peakVal 't_b_366+slope' baseVal
+ t_b_367 baseVal 't_b_367+slope' peakVal
+ t_b_368 peakVal 't_b_368+slope' baseVal
+ t_b_369 baseVal 't_b_369+slope' peakVal
+ t_b_370 peakVal 't_b_370+slope' baseVal
+ t_b_371 baseVal 't_b_371+slope' peakVal
+ t_b_372 peakVal 't_b_372+slope' baseVal
+ t_b_373 baseVal 't_b_373+slope' peakVal
+ t_b_374 peakVal 't_b_374+slope' baseVal
+ t_b_375 baseVal 't_b_375+slope' peakVal
+ t_b_376 peakVal 't_b_376+slope' baseVal
+ t_b_377 baseVal 't_b_377+slope' peakVal
+ t_b_378 peakVal 't_b_378+slope' baseVal
+ t_b_379 baseVal 't_b_379+slope' peakVal
+ t_b_380 peakVal 't_b_380+slope' baseVal
+ t_b_381 baseVal 't_b_381+slope' peakVal
+ t_b_382 peakVal 't_b_382+slope' baseVal
+ t_b_383 baseVal 't_b_383+slope' peakVal
+ t_b_384 peakVal 't_b_384+slope' baseVal
+ t_b_385 baseVal 't_b_385+slope' peakVal
+ t_b_386 peakVal 't_b_386+slope' baseVal
+ t_b_387 baseVal 't_b_387+slope' peakVal
+ t_b_388 peakVal 't_b_388+slope' baseVal
+ t_b_389 baseVal 't_b_389+slope' peakVal
+ t_b_390 peakVal 't_b_390+slope' baseVal
+ t_b_391 baseVal 't_b_391+slope' peakVal
+ t_b_392 peakVal 't_b_392+slope' baseVal
+ t_b_393 baseVal 't_b_393+slope' peakVal
+ t_b_394 peakVal 't_b_394+slope' baseVal
+ t_b_395 baseVal 't_b_395+slope' peakVal
+ t_b_396 peakVal 't_b_396+slope' baseVal
+ t_b_397 baseVal 't_b_397+slope' peakVal
+ t_b_398 peakVal 't_b_398+slope' baseVal
+ t_b_399 baseVal 't_b_399+slope' peakVal
+ t_b_400 peakVal 't_b_400+slope' baseVal
+ t_b_401 baseVal 't_b_401+slope' peakVal
+ t_b_402 peakVal 't_b_402+slope' baseVal
+ t_b_403 baseVal 't_b_403+slope' peakVal
+ t_b_404 peakVal 't_b_404+slope' baseVal
+ t_b_405 baseVal 't_b_405+slope' peakVal
+ t_b_406 peakVal 't_b_406+slope' baseVal
+ t_b_407 baseVal 't_b_407+slope' peakVal
+ t_b_408 peakVal 't_b_408+slope' baseVal
+ t_b_409 baseVal 't_b_409+slope' peakVal
+ t_b_410 peakVal 't_b_410+slope' baseVal
+ t_b_411 baseVal 't_b_411+slope' peakVal
+ t_b_412 peakVal 't_b_412+slope' baseVal
+ t_b_413 baseVal 't_b_413+slope' peakVal
+ t_b_414 peakVal 't_b_414+slope' baseVal
+ t_b_415 baseVal 't_b_415+slope' peakVal
+ t_b_416 peakVal 't_b_416+slope' baseVal
+ t_b_417 baseVal 't_b_417+slope' peakVal
+ t_b_418 peakVal 't_b_418+slope' baseVal
+ t_b_419 baseVal 't_b_419+slope' peakVal
+ t_b_420 peakVal 't_b_420+slope' baseVal
+ t_b_421 baseVal 't_b_421+slope' peakVal
+ t_b_422 peakVal 't_b_422+slope' baseVal
+ t_b_423 baseVal 't_b_423+slope' peakVal
+ t_b_424 peakVal 't_b_424+slope' baseVal
+ t_b_425 baseVal 't_b_425+slope' peakVal
+ t_b_426 peakVal 't_b_426+slope' baseVal
+ t_b_427 baseVal 't_b_427+slope' peakVal
+ t_b_428 peakVal 't_b_428+slope' baseVal
+ t_b_429 baseVal 't_b_429+slope' peakVal
+ t_b_430 peakVal 't_b_430+slope' baseVal
+ t_b_431 baseVal 't_b_431+slope' peakVal
+ t_b_432 peakVal 't_b_432+slope' baseVal
+ t_b_433 baseVal 't_b_433+slope' peakVal
+ t_b_434 peakVal 't_b_434+slope' baseVal
+ t_b_435 baseVal 't_b_435+slope' peakVal
+ t_b_436 peakVal 't_b_436+slope' baseVal
+ t_b_437 baseVal 't_b_437+slope' peakVal
+ t_b_438 peakVal 't_b_438+slope' baseVal
+ t_b_439 baseVal 't_b_439+slope' peakVal
+ t_b_440 peakVal 't_b_440+slope' baseVal
+ t_b_441 baseVal 't_b_441+slope' peakVal
+ t_b_442 peakVal 't_b_442+slope' baseVal
+ t_b_443 baseVal 't_b_443+slope' peakVal
+ t_b_444 peakVal 't_b_444+slope' baseVal
+ t_b_445 baseVal 't_b_445+slope' peakVal
+ t_b_446 peakVal 't_b_446+slope' baseVal
+ t_b_447 baseVal 't_b_447+slope' peakVal
+ t_b_448 peakVal 't_b_448+slope' baseVal
+ t_b_449 baseVal 't_b_449+slope' peakVal
+ t_b_450 peakVal 't_b_450+slope' baseVal
+ t_b_451 baseVal 't_b_451+slope' peakVal
+ t_b_452 peakVal 't_b_452+slope' baseVal
+ t_b_453 baseVal 't_b_453+slope' peakVal
+ t_b_454 peakVal 't_b_454+slope' baseVal
+ t_b_455 baseVal 't_b_455+slope' peakVal
+ t_b_456 peakVal 't_b_456+slope' baseVal
+ t_b_457 baseVal 't_b_457+slope' peakVal
+ t_b_458 peakVal 't_b_458+slope' baseVal
+ t_b_459 baseVal 't_b_459+slope' peakVal
+ t_b_460 peakVal 't_b_460+slope' baseVal
+ t_b_461 baseVal 't_b_461+slope' peakVal
+ t_b_462 peakVal 't_b_462+slope' baseVal
+ t_b_463 baseVal 't_b_463+slope' peakVal
+ t_b_464 peakVal 't_b_464+slope' baseVal
+ t_b_465 baseVal 't_b_465+slope' peakVal
+ t_b_466 peakVal 't_b_466+slope' baseVal
+ t_b_467 baseVal 't_b_467+slope' peakVal
+ t_b_468 peakVal 't_b_468+slope' baseVal
+ t_b_469 baseVal 't_b_469+slope' peakVal
+ t_b_470 peakVal 't_b_470+slope' baseVal
+ t_b_471 baseVal 't_b_471+slope' peakVal
+ t_b_472 peakVal 't_b_472+slope' baseVal
+ t_b_473 baseVal 't_b_473+slope' peakVal
+ t_b_474 peakVal 't_b_474+slope' baseVal
+ t_b_475 baseVal 't_b_475+slope' peakVal
+ t_b_476 peakVal 't_b_476+slope' baseVal
+ t_b_477 baseVal 't_b_477+slope' peakVal
+ t_b_478 peakVal 't_b_478+slope' baseVal
+ t_b_479 baseVal 't_b_479+slope' peakVal
+ t_b_480 peakVal 't_b_480+slope' baseVal
+ t_b_481 baseVal 't_b_481+slope' peakVal
+ t_b_482 peakVal 't_b_482+slope' baseVal
+ t_b_483 baseVal 't_b_483+slope' peakVal
+ t_b_484 peakVal 't_b_484+slope' baseVal
+ t_b_485 baseVal 't_b_485+slope' peakVal
+ t_b_486 peakVal 't_b_486+slope' baseVal
+ t_b_487 baseVal 't_b_487+slope' peakVal
+ t_b_488 peakVal 't_b_488+slope' baseVal
+ t_b_489 baseVal 't_b_489+slope' peakVal
+ t_b_490 peakVal 't_b_490+slope' baseVal
+ t_b_491 baseVal 't_b_491+slope' peakVal
+ t_b_492 peakVal 't_b_492+slope' baseVal
+ t_b_493 baseVal 't_b_493+slope' peakVal
+ t_b_494 peakVal 't_b_494+slope' baseVal
+ t_b_495 baseVal 't_b_495+slope' peakVal
+ t_b_496 peakVal 't_b_496+slope' baseVal
+ t_b_497 baseVal 't_b_497+slope' peakVal
+ t_b_498 peakVal 't_b_498+slope' baseVal
+ t_b_499 baseVal 't_b_499+slope' peakVal
+ t_b_500 peakVal 't_b_500+slope' baseVal
+ t_b_501 baseVal 't_b_501+slope' peakVal
+ t_b_502 peakVal 't_b_502+slope' baseVal
+ t_b_503 baseVal 't_b_503+slope' peakVal
+ t_b_504 peakVal 't_b_504+slope' baseVal
+ t_b_505 baseVal 't_b_505+slope' peakVal
+ t_b_506 peakVal 't_b_506+slope' baseVal
+ t_b_507 baseVal 't_b_507+slope' peakVal
+ t_b_508 peakVal 't_b_508+slope' baseVal
+ t_b_509 baseVal 't_b_509+slope' peakVal
+ t_b_510 peakVal 't_b_510+slope' baseVal
+ t_b_511 baseVal 't_b_511+slope' peakVal
+ t_b_512 peakVal 't_b_512+slope' baseVal
+ t_b_513 baseVal 't_b_513+slope' peakVal
+ t_b_514 peakVal 't_b_514+slope' baseVal
+ t_b_515 baseVal 't_b_515+slope' peakVal
+ t_b_516 peakVal 't_b_516+slope' baseVal
+ t_b_517 baseVal 't_b_517+slope' peakVal
+ t_b_518 peakVal 't_b_518+slope' baseVal
+ t_b_519 baseVal 't_b_519+slope' peakVal
+ t_b_520 peakVal 't_b_520+slope' baseVal
+ t_b_521 baseVal 't_b_521+slope' peakVal
+ t_b_522 peakVal 't_b_522+slope' baseVal
+ t_b_523 baseVal 't_b_523+slope' peakVal
+ t_b_524 peakVal 't_b_524+slope' baseVal
+ t_b_525 baseVal 't_b_525+slope' peakVal
+ t_b_526 peakVal 't_b_526+slope' baseVal
+ t_b_527 baseVal 't_b_527+slope' peakVal
+ t_b_528 peakVal 't_b_528+slope' baseVal
+ t_b_529 baseVal 't_b_529+slope' peakVal
+ t_b_530 peakVal 't_b_530+slope' baseVal
+ t_b_531 baseVal 't_b_531+slope' peakVal
+ t_b_532 peakVal 't_b_532+slope' baseVal
+ t_b_533 baseVal 't_b_533+slope' peakVal
+ t_b_534 peakVal 't_b_534+slope' baseVal
+ t_b_535 baseVal 't_b_535+slope' peakVal
+ t_b_536 peakVal 't_b_536+slope' baseVal
+ t_b_537 baseVal 't_b_537+slope' peakVal
+ t_b_538 peakVal 't_b_538+slope' baseVal
+ t_b_539 baseVal 't_b_539+slope' peakVal
+ t_b_540 peakVal 't_b_540+slope' baseVal
+ t_b_541 baseVal 't_b_541+slope' peakVal
+ t_b_542 peakVal 't_b_542+slope' baseVal
+ t_b_543 baseVal 't_b_543+slope' peakVal
+ t_b_544 peakVal 't_b_544+slope' baseVal
+ t_b_545 baseVal 't_b_545+slope' peakVal
+ t_b_546 peakVal 't_b_546+slope' baseVal
+ t_b_547 baseVal 't_b_547+slope' peakVal
+ t_b_548 peakVal 't_b_548+slope' baseVal
+ t_b_549 baseVal 't_b_549+slope' peakVal
+ t_b_550 peakVal 't_b_550+slope' baseVal
+ t_b_551 baseVal 't_b_551+slope' peakVal
+ t_b_552 peakVal 't_b_552+slope' baseVal
+ t_b_553 baseVal 't_b_553+slope' peakVal
+ t_b_554 peakVal 't_b_554+slope' baseVal
+ t_b_555 baseVal 't_b_555+slope' peakVal
+ t_b_556 peakVal 't_b_556+slope' baseVal
+ t_b_557 baseVal 't_b_557+slope' peakVal
+ t_b_558 peakVal 't_b_558+slope' baseVal
+ t_b_559 baseVal 't_b_559+slope' peakVal
+ t_b_560 peakVal 't_b_560+slope' baseVal
+ t_b_561 baseVal 't_b_561+slope' peakVal
+ t_b_562 peakVal 't_b_562+slope' baseVal
+ t_b_563 baseVal 't_b_563+slope' peakVal
+ t_b_564 peakVal 't_b_564+slope' baseVal
+ t_b_565 baseVal 't_b_565+slope' peakVal
+ t_b_566 peakVal 't_b_566+slope' baseVal
+ t_b_567 baseVal 't_b_567+slope' peakVal
+ t_b_568 peakVal 't_b_568+slope' baseVal
+ t_b_569 baseVal 't_b_569+slope' peakVal
+ t_b_570 peakVal 't_b_570+slope' baseVal
+ t_b_571 baseVal 't_b_571+slope' peakVal
+ t_b_572 peakVal 't_b_572+slope' baseVal
+ t_b_573 baseVal 't_b_573+slope' peakVal
+ t_b_574 peakVal 't_b_574+slope' baseVal
+ t_b_575 baseVal 't_b_575+slope' peakVal
+ t_b_576 peakVal 't_b_576+slope' baseVal
+ t_b_577 baseVal 't_b_577+slope' peakVal
+ t_b_578 peakVal 't_b_578+slope' baseVal
+ t_b_579 baseVal 't_b_579+slope' peakVal
+ t_b_580 peakVal 't_b_580+slope' baseVal
+ t_b_581 baseVal 't_b_581+slope' peakVal
+ t_b_582 peakVal 't_b_582+slope' baseVal
+ t_b_583 baseVal 't_b_583+slope' peakVal
+ t_b_584 peakVal 't_b_584+slope' baseVal
+ t_b_585 baseVal 't_b_585+slope' peakVal
+ t_b_586 peakVal 't_b_586+slope' baseVal
+ t_b_587 baseVal 't_b_587+slope' peakVal
+ t_b_588 peakVal 't_b_588+slope' baseVal
+ t_b_589 baseVal 't_b_589+slope' peakVal
+ t_b_590 peakVal 't_b_590+slope' baseVal
+ t_b_591 baseVal 't_b_591+slope' peakVal
+ t_b_592 peakVal 't_b_592+slope' baseVal
+ t_b_593 baseVal 't_b_593+slope' peakVal
+ t_b_594 peakVal 't_b_594+slope' baseVal
+ t_b_595 baseVal 't_b_595+slope' peakVal
+ t_b_596 peakVal 't_b_596+slope' baseVal
+ t_b_597 baseVal 't_b_597+slope' peakVal
+ t_b_598 peakVal 't_b_598+slope' baseVal
+ t_b_599 baseVal 't_b_599+slope' peakVal
+ t_b_600 peakVal 't_b_600+slope' baseVal
+ t_b_601 baseVal 't_b_601+slope' peakVal
+ t_b_602 peakVal 't_b_602+slope' baseVal
+ t_b_603 baseVal 't_b_603+slope' peakVal
+ t_b_604 peakVal 't_b_604+slope' baseVal
+ t_b_605 baseVal 't_b_605+slope' peakVal
+ t_b_606 peakVal 't_b_606+slope' baseVal
+ t_b_607 baseVal 't_b_607+slope' peakVal
+ t_b_608 peakVal 't_b_608+slope' baseVal
+ t_b_609 baseVal 't_b_609+slope' peakVal
+ t_b_610 peakVal 't_b_610+slope' baseVal
+ t_b_611 baseVal 't_b_611+slope' peakVal
+ t_b_612 peakVal 't_b_612+slope' baseVal
+ t_b_613 baseVal 't_b_613+slope' peakVal
+ t_b_614 peakVal 't_b_614+slope' baseVal
+ t_b_615 baseVal 't_b_615+slope' peakVal
+ t_b_616 peakVal 't_b_616+slope' baseVal
+ t_b_617 baseVal 't_b_617+slope' peakVal
+ t_b_618 peakVal 't_b_618+slope' baseVal
+ t_b_619 baseVal 't_b_619+slope' peakVal
+ t_b_620 peakVal 't_b_620+slope' baseVal
+ t_b_621 baseVal 't_b_621+slope' peakVal
+ t_b_622 peakVal 't_b_622+slope' baseVal
+ t_b_623 baseVal 't_b_623+slope' peakVal
+ t_b_624 peakVal 't_b_624+slope' baseVal
+ t_b_625 baseVal 't_b_625+slope' peakVal
+ t_b_626 peakVal 't_b_626+slope' baseVal
+ t_b_627 baseVal 't_b_627+slope' peakVal
+ t_b_628 peakVal 't_b_628+slope' baseVal
+ t_b_629 baseVal 't_b_629+slope' peakVal
+ t_b_630 peakVal 't_b_630+slope' baseVal
+ t_b_631 baseVal 't_b_631+slope' peakVal
+ t_b_632 peakVal 't_b_632+slope' baseVal
+ t_b_633 baseVal 't_b_633+slope' peakVal
+ t_b_634 peakVal 't_b_634+slope' baseVal
+ t_b_635 baseVal 't_b_635+slope' peakVal
+ t_b_636 peakVal 't_b_636+slope' baseVal
+ t_b_637 baseVal 't_b_637+slope' peakVal
+ t_b_638 peakVal 't_b_638+slope' baseVal
+ t_b_639 baseVal 't_b_639+slope' peakVal
+ t_b_640 peakVal 't_b_640+slope' baseVal
+ t_b_641 baseVal 't_b_641+slope' peakVal
+ t_b_642 peakVal 't_b_642+slope' baseVal
+ t_b_643 baseVal 't_b_643+slope' peakVal
+ t_b_644 peakVal 't_b_644+slope' baseVal
+ t_b_645 baseVal 't_b_645+slope' peakVal
+ t_b_646 peakVal 't_b_646+slope' baseVal
+ t_b_647 baseVal 't_b_647+slope' peakVal
+ t_b_648 peakVal 't_b_648+slope' baseVal
+ t_b_649 baseVal 't_b_649+slope' peakVal
+ t_b_650 peakVal 't_b_650+slope' baseVal
+ t_b_651 baseVal 't_b_651+slope' peakVal
+ t_b_652 peakVal 't_b_652+slope' baseVal
+ t_b_653 baseVal 't_b_653+slope' peakVal
+ t_b_654 peakVal 't_b_654+slope' baseVal
+ t_b_655 baseVal 't_b_655+slope' peakVal
+ t_b_656 peakVal 't_b_656+slope' baseVal
+ t_b_657 baseVal 't_b_657+slope' peakVal
+ t_b_658 peakVal 't_b_658+slope' baseVal
+ t_b_659 baseVal 't_b_659+slope' peakVal
+ t_b_660 peakVal 't_b_660+slope' baseVal
+ t_b_661 baseVal 't_b_661+slope' peakVal
+ t_b_662 peakVal 't_b_662+slope' baseVal
+ t_b_663 baseVal 't_b_663+slope' peakVal
+ t_b_664 peakVal 't_b_664+slope' baseVal
+ t_b_665 baseVal 't_b_665+slope' peakVal
+ t_b_666 peakVal 't_b_666+slope' baseVal
+ t_b_667 baseVal 't_b_667+slope' peakVal
+ t_b_668 peakVal 't_b_668+slope' baseVal
+ t_b_669 baseVal 't_b_669+slope' peakVal
+ t_b_670 peakVal 't_b_670+slope' baseVal
+ t_b_671 baseVal 't_b_671+slope' peakVal
+ t_b_672 peakVal 't_b_672+slope' baseVal
+ t_b_673 baseVal 't_b_673+slope' peakVal
+ t_b_674 peakVal 't_b_674+slope' baseVal
+ t_b_675 baseVal 't_b_675+slope' peakVal
+ t_b_676 peakVal 't_b_676+slope' baseVal
+ t_b_677 baseVal 't_b_677+slope' peakVal
+ t_b_678 peakVal 't_b_678+slope' baseVal
+ t_b_679 baseVal 't_b_679+slope' peakVal
+ t_b_680 peakVal 't_b_680+slope' baseVal
+ t_b_681 baseVal 't_b_681+slope' peakVal
+ t_b_682 peakVal 't_b_682+slope' baseVal
+ t_b_683 baseVal 't_b_683+slope' peakVal
+ t_b_684 peakVal 't_b_684+slope' baseVal
+ t_b_685 baseVal 't_b_685+slope' peakVal
+ t_b_686 peakVal 't_b_686+slope' baseVal
+ t_b_687 baseVal 't_b_687+slope' peakVal
+ t_b_688 peakVal 't_b_688+slope' baseVal
+ t_b_689 baseVal 't_b_689+slope' peakVal
+ t_b_690 peakVal 't_b_690+slope' baseVal
+ t_b_691 baseVal 't_b_691+slope' peakVal
+ t_b_692 peakVal 't_b_692+slope' baseVal
+ t_b_693 baseVal 't_b_693+slope' peakVal
+ t_b_694 peakVal 't_b_694+slope' baseVal
+ t_b_695 baseVal 't_b_695+slope' peakVal
+ t_b_696 peakVal 't_b_696+slope' baseVal
+ t_b_697 baseVal 't_b_697+slope' peakVal
+ t_b_698 peakVal 't_b_698+slope' baseVal
+ t_b_699 baseVal 't_b_699+slope' peakVal
+ t_b_700 peakVal 't_b_700+slope' baseVal
+ t_b_701 baseVal 't_b_701+slope' peakVal
+ t_b_702 peakVal 't_b_702+slope' baseVal
+ t_b_703 baseVal 't_b_703+slope' peakVal
+ t_b_704 peakVal 't_b_704+slope' baseVal
+ t_b_705 baseVal 't_b_705+slope' peakVal
+ t_b_706 peakVal 't_b_706+slope' baseVal
+ t_b_707 baseVal 't_b_707+slope' peakVal
+ t_b_708 peakVal 't_b_708+slope' baseVal
+ t_b_709 baseVal 't_b_709+slope' peakVal
+ t_b_710 peakVal 't_b_710+slope' baseVal
+ t_b_711 baseVal 't_b_711+slope' peakVal
+ t_b_712 peakVal 't_b_712+slope' baseVal
+ t_b_713 baseVal 't_b_713+slope' peakVal
+ t_b_714 peakVal 't_b_714+slope' baseVal
+ t_b_715 baseVal 't_b_715+slope' peakVal
+ t_b_716 peakVal 't_b_716+slope' baseVal
+ t_b_717 baseVal 't_b_717+slope' peakVal
+ t_b_718 peakVal 't_b_718+slope' baseVal
+ t_b_719 baseVal 't_b_719+slope' peakVal
+ t_b_720 peakVal 't_b_720+slope' baseVal
+ t_b_721 baseVal 't_b_721+slope' peakVal
+ t_b_722 peakVal 't_b_722+slope' baseVal
+ t_b_723 baseVal 't_b_723+slope' peakVal
+ t_b_724 peakVal 't_b_724+slope' baseVal
+ t_b_725 baseVal 't_b_725+slope' peakVal
+ t_b_726 peakVal 't_b_726+slope' baseVal
+ t_b_727 baseVal 't_b_727+slope' peakVal
+ t_b_728 peakVal 't_b_728+slope' baseVal
+ t_b_729 baseVal 't_b_729+slope' peakVal
+ t_b_730 peakVal 't_b_730+slope' baseVal
+ t_b_731 baseVal 't_b_731+slope' peakVal
+ t_b_732 peakVal 't_b_732+slope' baseVal
+ t_b_733 baseVal 't_b_733+slope' peakVal
+ t_b_734 peakVal 't_b_734+slope' baseVal
+ t_b_735 baseVal 't_b_735+slope' peakVal
+ t_b_736 peakVal 't_b_736+slope' baseVal
+ t_b_737 baseVal 't_b_737+slope' peakVal
+ t_b_738 peakVal 't_b_738+slope' baseVal
+ t_b_739 baseVal 't_b_739+slope' peakVal
+ t_b_740 peakVal 't_b_740+slope' baseVal
+ t_b_741 baseVal 't_b_741+slope' peakVal
+ t_b_742 peakVal 't_b_742+slope' baseVal
+ t_b_743 baseVal 't_b_743+slope' peakVal
+ t_b_744 peakVal 't_b_744+slope' baseVal
+ t_b_745 baseVal 't_b_745+slope' peakVal
+ t_b_746 peakVal 't_b_746+slope' baseVal
+ t_b_747 baseVal 't_b_747+slope' peakVal
+ t_b_748 peakVal 't_b_748+slope' baseVal
+ t_b_749 baseVal 't_b_749+slope' peakVal
+ t_b_750 peakVal 't_b_750+slope' baseVal
+ t_b_751 baseVal 't_b_751+slope' peakVal
+ t_b_752 peakVal 't_b_752+slope' baseVal
+ t_b_753 baseVal 't_b_753+slope' peakVal
+ t_b_754 peakVal 't_b_754+slope' baseVal
+ t_b_755 baseVal 't_b_755+slope' peakVal
+ t_b_756 peakVal 't_b_756+slope' baseVal
+ t_b_757 baseVal 't_b_757+slope' peakVal
+ t_b_758 peakVal 't_b_758+slope' baseVal
+ t_b_759 baseVal 't_b_759+slope' peakVal
+ t_b_760 peakVal 't_b_760+slope' baseVal
+ t_b_761 baseVal 't_b_761+slope' peakVal
+ t_b_762 peakVal 't_b_762+slope' baseVal
+ t_b_763 baseVal 't_b_763+slope' peakVal
+ t_b_764 peakVal 't_b_764+slope' baseVal
+ t_b_765 baseVal 't_b_765+slope' peakVal
+ t_b_766 peakVal 't_b_766+slope' baseVal
+ t_b_767 baseVal 't_b_767+slope' peakVal
+ t_b_768 peakVal 't_b_768+slope' baseVal
+ t_b_769 baseVal 't_b_769+slope' peakVal
+ t_b_770 peakVal 't_b_770+slope' baseVal
+ t_b_771 baseVal 't_b_771+slope' peakVal
+ t_b_772 peakVal 't_b_772+slope' baseVal
+ t_b_773 baseVal 't_b_773+slope' peakVal
+ t_b_774 peakVal 't_b_774+slope' baseVal
+ t_b_775 baseVal 't_b_775+slope' peakVal
+ t_b_776 peakVal 't_b_776+slope' baseVal
+ t_b_777 baseVal 't_b_777+slope' peakVal
+ t_b_778 peakVal 't_b_778+slope' baseVal
+ t_b_779 baseVal 't_b_779+slope' peakVal
+ t_b_780 peakVal 't_b_780+slope' baseVal
+ t_b_781 baseVal 't_b_781+slope' peakVal
+ t_b_782 peakVal 't_b_782+slope' baseVal
+ t_b_783 baseVal 't_b_783+slope' peakVal
+ t_b_784 peakVal 't_b_784+slope' baseVal
+ t_b_785 baseVal 't_b_785+slope' peakVal
+ t_b_786 peakVal 't_b_786+slope' baseVal
+ t_b_787 baseVal 't_b_787+slope' peakVal
+ t_b_788 peakVal 't_b_788+slope' baseVal
+ t_b_789 baseVal 't_b_789+slope' peakVal
+ t_b_790 peakVal 't_b_790+slope' baseVal
+ t_b_791 baseVal 't_b_791+slope' peakVal
+ t_b_792 peakVal 't_b_792+slope' baseVal
+ t_b_793 baseVal 't_b_793+slope' peakVal
+ t_b_794 peakVal 't_b_794+slope' baseVal
+ t_b_795 baseVal 't_b_795+slope' peakVal
+ t_b_796 peakVal 't_b_796+slope' baseVal
+ t_b_797 baseVal 't_b_797+slope' peakVal
+ t_b_798 peakVal 't_b_798+slope' baseVal
+ t_b_799 baseVal 't_b_799+slope' peakVal


*circuit

XBUFFER_A Input_A A VDD VDD GND GND BUF_X8
XBUFFER_B Input_B B VDD VDD GND GND BUF_X8
XCGATE A B Z VDD VDD GND GND CGATE
XBUFFER_Z Z Output VDD VDD GND GND BUF_X8
C_TERM Output GND 0.0779pF

.PROBE TRAN V(A) V(B) V(Z)
.TRAN 0.1ps tend
.END
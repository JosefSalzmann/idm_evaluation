* circuit: nor inv chain
simulator lang=spice

*.PARAM pw=<sed>pw<sed>as
.PARAM supp=0.8V slope=0.1fs
.PARAM t_init0=0.1ns t_init1=0.174ns
.PARAM baseVal=0V peakVal=0.8V tend=1.0ns


.LIB /home/s11777724/involution_tool_library_files/backend/spice/fet.inc CMG

* main circuit
.INCLUDE /home/s11777724/involution_tool_library_files/backend/spice/cell/NOR2_X1.sp

**** SPECTRE Back Annotation
.option spef='../place_and_route/generic_parasitics.spef'
****

.TEMP 25
.OPTION
+ INGOLD=2
+ PARHIER=LOCAL
*+ POST=CSDF
+ PROBE
+ BRIEF
+ ACCURATE
+ ABSVAR=0.0001
+ DVDT=2
+ RELTOL=1e-11
*+ DELMAX=100fs
+ dc_pivot_check=yes

* vdd
VDD VDD GND 0.8v

VIN IN_A GND PWL 0ns baseVal t_init0 baseVal 't_init0+slope' peakVal t_init1 peakVal 't_init1+slope' baseVal
VIN IN_B GND PWL 0ns baseVal t_init0 baseVal 't_init0+slope' peakVal t_init1 peakVal 't_init1+slope' baseVal

* circuit under test
X_NOR_STAGE_0_1 IN_A IN_B  STAGE_0_OUT_1 VDD VDD GND GND NOR2_X2
X_NOR_STAGE_0_2 IN_A IN_B  STAGE_0_OUT_2 VDD VDD GND GND NOR2_X2

X_NOR_STAGE_1_1 STAGE_0_OUT_1 STAGE_0_OUT_2  STAGE_1_OUT_1 VDD VDD GND GND NOR2_X2
X_NOR_STAGE_1_2 STAGE_0_OUT_1 STAGE_0_OUT_2  STAGE_1_OUT_2 VDD VDD GND GND NOR2_X2

X_NOR_STAGE_2_1 STAGE_1_OUT_1 STAGE_1_OUT_2  STAGE_2_OUT_1 VDD VDD GND GND NOR2_X2
X_NOR_STAGE_2_2 STAGE_1_OUT_1 STAGE_1_OUT_2  STAGE_2_OUT_2 VDD VDD GND GND NOR2_X2

X_NOR_STAGE_3_1 STAGE_2_OUT_1 STAGE_2_OUT_2  STAGE_3_OUT_1 VDD VDD GND GND NOR2_X2
X_NOR_STAGE_3_2 STAGE_2_OUT_1 STAGE_2_OUT_2  STAGE_3_OUT_2 VDD VDD GND GND NOR2_X2

X_NOR_STAGE_4_1 STAGE_3_OUT_1 STAGE_3_OUT_2  STAGE_4_OUT_1 VDD VDD GND GND NOR2_X2
X_NOR_STAGE_4_2 STAGE_3_OUT_1 STAGE_3_OUT_2  STAGE_4_OUT_2 VDD VDD GND GND NOR2_X2

X_NOR_STAGE_5_1 STAGE_4_OUT_1 STAGE_4_OUT_2  STAGE_5_OUT_1 VDD VDD GND GND NOR2_X2
X_NOR_STAGE_5_2 STAGE_4_OUT_1 STAGE_4_OUT_2  STAGE_5_OUT_2 VDD VDD GND GND NOR2_X2

X_NOR_STAGE_6_1 STAGE_5_OUT_1 STAGE_5_OUT_2  STAGE_6_OUT_1 VDD VDD GND GND NOR2_X2
X_NOR_STAGE_6_2 STAGE_5_OUT_1 STAGE_5_OUT_2  STAGE_6_OUT_2 VDD VDD GND GND NOR2_X2

X_NOR_STAGE_7_1 STAGE_6_OUT_1 STAGE_6_OUT_2  STAGE_7_OUT_1 VDD VDD GND GND NOR2_X2
X_NOR_STAGE_7_2 STAGE_6_OUT_1 STAGE_6_OUT_2  STAGE_7_OUT_2 VDD VDD GND GND NOR2_X2

X_NOR_STAGE_8_1 STAGE_7_OUT_1 STAGE_7_OUT_2  STAGE_8_OUT_1 VDD VDD GND GND NOR2_X2
X_NOR_STAGE_8_2 STAGE_7_OUT_1 STAGE_7_OUT_2  STAGE_8_OUT_2 VDD VDD GND GND NOR2_X2

X_NOR_STAGE_9_1 STAGE_8_OUT_1 STAGE_8_OUT_2  STAGE_9_OUT_1 VDD VDD GND GND NOR2_X2
X_NOR_STAGE_9_2 STAGE_8_OUT_1 STAGE_8_OUT_2  STAGE_9_OUT_2 VDD VDD GND GND NOR2_X2

X_NOR_STAGE_10_1 STAGE_9_OUT_1 STAGE_9_OUT_2  STAGE_10_OUT_1 VDD VDD GND GND NOR2_X2
X_NOR_STAGE_10_2 STAGE_9_OUT_1 STAGE_9_OUT_2  STAGE_10_OUT_2 VDD VDD GND GND NOR2_X2

X_NOR_STAGE_11_1 STAGE_10_OUT_1 STAGE_10_OUT_2  STAGE_11_OUT_1 VDD VDD GND GND NOR2_X2
X_NOR_STAGE_11_2 STAGE_10_OUT_1 STAGE_10_OUT_2  STAGE_11_OUT_2 VDD VDD GND GND NOR2_X2

X_NOR_STAGE_12_1 STAGE_11_OUT_1 STAGE_11_OUT_2  STAGE_12_OUT_1 VDD VDD GND GND NOR2_X2
X_NOR_STAGE_12_2 STAGE_11_OUT_1 STAGE_11_OUT_2  STAGE_12_OUT_2 VDD VDD GND GND NOR2_X2

X_NOR_STAGE_13_1 STAGE_12_OUT_1 STAGE_12_OUT_2  STAGE_13_OUT_1 VDD VDD GND GND NOR2_X2
X_NOR_STAGE_13_2 STAGE_12_OUT_1 STAGE_12_OUT_2  STAGE_13_OUT_2 VDD VDD GND GND NOR2_X2

X_NOR_STAGE_14_1 STAGE_13_OUT_1 STAGE_13_OUT_2  STAGE_14_OUT_1 VDD VDD GND GND NOR2_X2
X_NOR_STAGE_14_2 STAGE_13_OUT_1 STAGE_13_OUT_2  STAGE_14_OUT_2 VDD VDD GND GND NOR2_X2

X_NOR_STAGE_15_1 STAGE_14_OUT_1 STAGE_14_OUT_2  STAGE_15_OUT_1 VDD VDD GND GND NOR2_X2
X_NOR_STAGE_15_2 STAGE_14_OUT_1 STAGE_14_OUT_2  STAGE_15_OUT_2 VDD VDD GND GND NOR2_X2

X_NOR_STAGE_16_1 STAGE_15_OUT_1 STAGE_15_OUT_2  STAGE_16_OUT_1 VDD VDD GND GND NOR2_X2
X_NOR_STAGE_16_2 STAGE_15_OUT_1 STAGE_15_OUT_2  STAGE_16_OUT_2 VDD VDD GND GND NOR2_X2

X_NOR_STAGE_17_1 STAGE_16_OUT_1 STAGE_16_OUT_2  STAGE_17_OUT_1 VDD VDD GND GND NOR2_X2
X_NOR_STAGE_17_2 STAGE_16_OUT_1 STAGE_16_OUT_2  STAGE_17_OUT_2 VDD VDD GND GND NOR2_X2

X_NOR_STAGE_18_1 STAGE_17_OUT_1 STAGE_17_OUT_2  STAGE_18_OUT_1 VDD VDD GND GND NOR2_X2
X_NOR_STAGE_18_2 STAGE_17_OUT_1 STAGE_17_OUT_2  STAGE_18_OUT_2 VDD VDD GND GND NOR2_X2

X_NOR_STAGE_19_1 STAGE_18_OUT_1 STAGE_18_OUT_2  STAGE_19_OUT_1 VDD VDD GND GND NOR2_X2
X_NOR_STAGE_19_2 STAGE_18_OUT_1 STAGE_18_OUT_2  STAGE_19_OUT_2 VDD VDD GND GND NOR2_X2

X_NOR_STAGE_20_1 STAGE_19_OUT_1 STAGE_19_OUT_2  STAGE_20_OUT_1 VDD VDD GND GND NOR2_X2
X_NOR_STAGE_20_2 STAGE_19_OUT_1 STAGE_19_OUT_2  STAGE_20_OUT_2 VDD VDD GND GND NOR2_X2

X_NOR_STAGE_21_1 STAGE_20_OUT_1 STAGE_20_OUT_2  STAGE_21_OUT_1 VDD VDD GND GND NOR2_X2
X_NOR_STAGE_21_2 STAGE_20_OUT_1 STAGE_20_OUT_2  STAGE_21_OUT_2 VDD VDD GND GND NOR2_X2

X_NOR_STAGE_22_1 STAGE_21_OUT_1 STAGE_21_OUT_2  STAGE_22_OUT_1 VDD VDD GND GND NOR2_X2
X_NOR_STAGE_22_2 STAGE_21_OUT_1 STAGE_21_OUT_2  STAGE_22_OUT_2 VDD VDD GND GND NOR2_X2

X_NOR_STAGE_23_1 STAGE_22_OUT_1 STAGE_22_OUT_2  STAGE_23_OUT_1 VDD VDD GND GND NOR2_X2
X_NOR_STAGE_23_2 STAGE_22_OUT_1 STAGE_22_OUT_2  STAGE_23_OUT_2 VDD VDD GND GND NOR2_X2

X_NOR_STAGE_24_1 STAGE_23_OUT_1 STAGE_23_OUT_2  STAGE_24_OUT_1 VDD VDD GND GND NOR2_X2
X_NOR_STAGE_24_2 STAGE_23_OUT_1 STAGE_23_OUT_2  STAGE_24_OUT_2 VDD VDD GND GND NOR2_X2

X_NOR_STAGE_25_1 STAGE_24_OUT_1 STAGE_24_OUT_2  STAGE_25_OUT_1 VDD VDD GND GND NOR2_X2
X_NOR_STAGE_25_2 STAGE_24_OUT_1 STAGE_24_OUT_2  STAGE_25_OUT_2 VDD VDD GND GND NOR2_X2

X_NOR_STAGE_26_1 STAGE_25_OUT_1 STAGE_25_OUT_2  STAGE_26_OUT_1 VDD VDD GND GND NOR2_X2
X_NOR_STAGE_26_2 STAGE_25_OUT_1 STAGE_25_OUT_2  STAGE_26_OUT_2 VDD VDD GND GND NOR2_X2

X_NOR_STAGE_27_1 STAGE_26_OUT_1 STAGE_26_OUT_2  STAGE_27_OUT_1 VDD VDD GND GND NOR2_X2
X_NOR_STAGE_27_2 STAGE_26_OUT_1 STAGE_26_OUT_2  STAGE_27_OUT_2 VDD VDD GND GND NOR2_X2

X_NOR_STAGE_28_1 STAGE_27_OUT_1 STAGE_27_OUT_2  STAGE_28_OUT_1 VDD VDD GND GND NOR2_X2
X_NOR_STAGE_28_2 STAGE_27_OUT_1 STAGE_27_OUT_2  STAGE_28_OUT_2 VDD VDD GND GND NOR2_X2

X_NOR_STAGE_29_1 STAGE_28_OUT_1 STAGE_28_OUT_2  STAGE_29_OUT_1 VDD VDD GND GND NOR2_X2
X_NOR_STAGE_29_2 STAGE_28_OUT_1 STAGE_28_OUT_2  STAGE_29_OUT_2 VDD VDD GND GND NOR2_X2

X_NOR_STAGE_30_1 STAGE_29_OUT_1 STAGE_29_OUT_2  STAGE_30_OUT_1 VDD VDD GND GND NOR2_X2
X_NOR_STAGE_30_2 STAGE_29_OUT_1 STAGE_29_OUT_2  STAGE_30_OUT_2 VDD VDD GND GND NOR2_X2

X_NOR_STAGE_31_1 STAGE_30_OUT_1 STAGE_30_OUT_2  STAGE_31_OUT_1 VDD VDD GND GND NOR2_X2
X_NOR_STAGE_31_2 STAGE_30_OUT_1 STAGE_30_OUT_2  STAGE_31_OUT_2 VDD VDD GND GND NOR2_X2

X_NOR_STAGE_32_1 STAGE_31_OUT_1 STAGE_31_OUT_2  STAGE_32_OUT_1 VDD VDD GND GND NOR2_X2
X_NOR_STAGE_32_2 STAGE_31_OUT_1 STAGE_31_OUT_2  STAGE_32_OUT_2 VDD VDD GND GND NOR2_X2

X_NOR_STAGE_33_1 STAGE_32_OUT_1 STAGE_32_OUT_2  STAGE_33_OUT_1 VDD VDD GND GND NOR2_X2
X_NOR_STAGE_33_2 STAGE_32_OUT_1 STAGE_32_OUT_2  STAGE_33_OUT_2 VDD VDD GND GND NOR2_X2

X_NOR_STAGE_34_1 STAGE_33_OUT_1 STAGE_33_OUT_2  STAGE_34_OUT_1 VDD VDD GND GND NOR2_X2
X_NOR_STAGE_34_2 STAGE_33_OUT_1 STAGE_33_OUT_2  STAGE_34_OUT_2 VDD VDD GND GND NOR2_X2

X_NOR_STAGE_35_1 STAGE_34_OUT_1 STAGE_34_OUT_2  STAGE_35_OUT_1 VDD VDD GND GND NOR2_X2
X_NOR_STAGE_35_2 STAGE_34_OUT_1 STAGE_34_OUT_2  STAGE_35_OUT_2 VDD VDD GND GND NOR2_X2

X_NOR_STAGE_36_1 STAGE_35_OUT_1 STAGE_35_OUT_2  STAGE_36_OUT_1 VDD VDD GND GND NOR2_X2
X_NOR_STAGE_36_2 STAGE_35_OUT_1 STAGE_35_OUT_2  STAGE_36_OUT_2 VDD VDD GND GND NOR2_X2

X_NOR_STAGE_37_1 STAGE_36_OUT_1 STAGE_36_OUT_2  STAGE_37_OUT_1 VDD VDD GND GND NOR2_X2
X_NOR_STAGE_37_2 STAGE_36_OUT_1 STAGE_36_OUT_2  STAGE_37_OUT_2 VDD VDD GND GND NOR2_X2

X_NOR_STAGE_38_1 STAGE_37_OUT_1 STAGE_37_OUT_2  STAGE_38_OUT_1 VDD VDD GND GND NOR2_X2
X_NOR_STAGE_38_2 STAGE_37_OUT_1 STAGE_37_OUT_2  STAGE_38_OUT_2 VDD VDD GND GND NOR2_X2

X_NOR_STAGE_39_1 STAGE_38_OUT_1 STAGE_38_OUT_2  STAGE_39_OUT_1 VDD VDD GND GND NOR2_X2
X_NOR_STAGE_39_2 STAGE_38_OUT_1 STAGE_38_OUT_2  STAGE_39_OUT_2 VDD VDD GND GND NOR2_X2

X_NOR_STAGE_40_1 STAGE_39_OUT_1 STAGE_39_OUT_2  STAGE_40_OUT_1 VDD VDD GND GND NOR2_X2
X_NOR_STAGE_40_2 STAGE_39_OUT_1 STAGE_39_OUT_2  STAGE_40_OUT_2 VDD VDD GND GND NOR2_X2

X_NOR_STAGE_41_1 STAGE_40_OUT_1 STAGE_40_OUT_2  STAGE_41_OUT_1 VDD VDD GND GND NOR2_X2
X_NOR_STAGE_41_2 STAGE_40_OUT_1 STAGE_40_OUT_2  STAGE_41_OUT_2 VDD VDD GND GND NOR2_X2

X_NOR_STAGE_42_1 STAGE_41_OUT_1 STAGE_41_OUT_2  STAGE_42_OUT_1 VDD VDD GND GND NOR2_X2
X_NOR_STAGE_42_2 STAGE_41_OUT_1 STAGE_41_OUT_2  STAGE_42_OUT_2 VDD VDD GND GND NOR2_X2

X_NOR_STAGE_43_1 STAGE_42_OUT_1 STAGE_42_OUT_2  STAGE_43_OUT_1 VDD VDD GND GND NOR2_X2
X_NOR_STAGE_43_2 STAGE_42_OUT_1 STAGE_42_OUT_2  STAGE_43_OUT_2 VDD VDD GND GND NOR2_X2

X_NOR_STAGE_44_1 STAGE_43_OUT_1 STAGE_43_OUT_2  STAGE_44_OUT_1 VDD VDD GND GND NOR2_X2
X_NOR_STAGE_44_2 STAGE_43_OUT_1 STAGE_43_OUT_2  STAGE_44_OUT_2 VDD VDD GND GND NOR2_X2

X_NOR_STAGE_45_1 STAGE_44_OUT_1 STAGE_44_OUT_2  STAGE_45_OUT_1 VDD VDD GND GND NOR2_X2
X_NOR_STAGE_45_2 STAGE_44_OUT_1 STAGE_44_OUT_2  STAGE_45_OUT_2 VDD VDD GND GND NOR2_X2

X_NOR_STAGE_46_1 STAGE_45_OUT_1 STAGE_45_OUT_2  STAGE_46_OUT_1 VDD VDD GND GND NOR2_X2
X_NOR_STAGE_46_2 STAGE_45_OUT_1 STAGE_45_OUT_2  STAGE_46_OUT_2 VDD VDD GND GND NOR2_X2

X_NOR_STAGE_47_1 STAGE_46_OUT_1 STAGE_46_OUT_2  STAGE_47_OUT_1 VDD VDD GND GND NOR2_X2
X_NOR_STAGE_47_2 STAGE_46_OUT_1 STAGE_46_OUT_2  STAGE_47_OUT_2 VDD VDD GND GND NOR2_X2

X_NOR_STAGE_48_1 STAGE_47_OUT_1 STAGE_47_OUT_2  STAGE_48_OUT_1 VDD VDD GND GND NOR2_X2
X_NOR_STAGE_48_2 STAGE_47_OUT_1 STAGE_47_OUT_2  STAGE_48_OUT_2 VDD VDD GND GND NOR2_X2

X_NOR_STAGE_49_1 STAGE_48_OUT_1 STAGE_48_OUT_2  STAGE_49_OUT_1 VDD VDD GND GND NOR2_X2
X_NOR_STAGE_49_2 STAGE_48_OUT_1 STAGE_48_OUT_2  STAGE_49_OUT_2 VDD VDD GND GND NOR2_X2

X_NOR_STAGE_50_1 STAGE_49_OUT_1 STAGE_49_OUT_2  STAGE_50_OUT_1 VDD VDD GND GND NOR2_X2
X_NOR_STAGE_50_2 STAGE_49_OUT_1 STAGE_49_OUT_2  STAGE_50_OUT_2 VDD VDD GND GND NOR2_X2

X_NOR_STAGE_51_1 STAGE_50_OUT_1 STAGE_50_OUT_2  STAGE_51_OUT_1 VDD VDD GND GND NOR2_X2
X_NOR_STAGE_51_2 STAGE_50_OUT_1 STAGE_50_OUT_2  STAGE_51_OUT_2 VDD VDD GND GND NOR2_X2

X_NOR_STAGE_52_1 STAGE_51_OUT_1 STAGE_51_OUT_2  STAGE_52_OUT_1 VDD VDD GND GND NOR2_X2
X_NOR_STAGE_52_2 STAGE_51_OUT_1 STAGE_51_OUT_2  STAGE_52_OUT_2 VDD VDD GND GND NOR2_X2

X_NOR_STAGE_53_1 STAGE_52_OUT_1 STAGE_52_OUT_2  STAGE_53_OUT_1 VDD VDD GND GND NOR2_X2
X_NOR_STAGE_53_2 STAGE_52_OUT_1 STAGE_52_OUT_2  STAGE_53_OUT_2 VDD VDD GND GND NOR2_X2

C_STAGE_53_TERM_1 STAGE_53_OUT_1 GND 0.01PF
C_STAGE_53_TERM_2 STAGE_53_OUT_2 GND 0.01PF
C_TERM myout GND 0.0779pF

.PROBE TRAN V(myin) V(STAGE1) V(STAGE2) V(STAGE3) V(STAGE4) V(STAGE5) V(STAGE6) V(STAGE7) V(STAGE8) V(STAGE9) V(STAGE10) V(STAGE11) V(STAGE12) V(STAGE13) V(STAGE14) V(STAGE15) V(STAGE16) V(STAGE17) V(STAGE18) V(STAGE19) V(STAGE20) V(STAGE21) V(STAGE22) V(STAGE23) V(STAGE24) V(STAGE25) V(STAGE26) V(STAGE27) V(STAGE28) V(STAGE29) V(STAGE30) V(STAGE31) V(STAGE32) V(STAGE33) V(STAGE34) V(STAGE35) V(STAGE36) V(STAGE37) V(STAGE38) V(STAGE39) V(STAGE40) V(STAGE41) V(STAGE42) V(STAGE43) V(STAGE44) V(STAGE45) V(STAGE46) V(STAGE47) V(STAGE48) V(STAGE49) V(STAGE50) V(STAGE51) V(STAGE52) V(STAGE53) V(STAGE54) V(STAGE55) V(STAGE56) V(STAGE57) V(STAGE58) V(STAGE59) V(STAGE60) V(STAGE61) V(STAGE62) V(STAGE63) V(STAGE64) V(STAGE65) V(STAGE66) V(STAGE67) V(STAGE68) V(STAGE69) V(STAGE70) V(STAGE71) V(STAGE72) V(STAGE73) V(STAGE74) V(STAGE75) V(STAGE76) V(STAGE77) V(STAGE78) V(STAGE79) V(STAGE80) V(STAGE81) V(STAGE82) V(STAGE83) V(STAGE84) V(STAGE85) V(STAGE86) V(STAGE87) V(STAGE88) V(STAGE89) V(STAGE90) V(STAGE91) V(STAGE92) V(STAGE93) V(STAGE94) V(STAGE95) V(STAGE96) V(STAGE97) V(STAGE98) V(STAGE99) V(STAGE100) V(STAGE101) V(STAGE102) V(STAGE103) V(STAGE104) V(STAGE105) V(STAGE106) V(STAGE107) V(STAGE108) V(STAGE109) V(STAGE110) V(STAGE111) V(STAGE112) V(STAGE113) V(STAGE114) V(STAGE115)
.TRAN 0.1ps tend
.END

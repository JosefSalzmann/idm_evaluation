module c880_NOR_template (N1_PWL,N8_PWL,N13_PWL,N17_PWL,N26_PWL,N29_PWL,N36_PWL,N42_PWL,N51_PWL,N55_PWL,
            N59_PWL,N68_PWL,N72_PWL,N73_PWL,N74_PWL,N75_PWL,N80_PWL,N85_PWL,N86_PWL,N87_PWL,
            N88_PWL,N89_PWL,N90_PWL,N91_PWL,N96_PWL,N101_PWL,N106_PWL,N111_PWL,N116_PWL,N121_PWL,
            N126_PWL,N130_PWL,N135_PWL,N138_PWL,N143_PWL,N146_PWL,N149_PWL,N152_PWL,N153_PWL,N156_PWL,
            N159_PWL,N165_PWL,N171_PWL,N177_PWL,N183_PWL,N189_PWL,N195_PWL,N201_PWL,N207_PWL,N210_PWL,
            N219_PWL,N228_PWL,N237_PWL,N246_PWL,N255_PWL,N259_PWL,N260_PWL,N261_PWL,N267_PWL,N268_PWL,
            N388_TERMINATION,N389_TERMINATION,N390_TERMINATION,N391_TERMINATION,N418_TERMINATION,
            N419_TERMINATION,N420_TERMINATION,N421_TERMINATION,N422_TERMINATION,N423_TERMINATION,
            N446_TERMINATION,N447_TERMINATION,N448_TERMINATION,N449_TERMINATION,N450_TERMINATION,
            N767_TERMINATION,N768_TERMINATION,N850_TERMINATION,N863_TERMINATION,N864_TERMINATION,
            N865_TERMINATION,N866_TERMINATION,N874_TERMINATION,N878_TERMINATION,N879_TERMINATION,
            N880_TERMINATION);

      input N1_PWL,N8_PWL,N13_PWL,N17_PWL,N26_PWL,N29_PWL,N36_PWL,N42_PWL,N51_PWL,N55_PWL,
            N59_PWL,N68_PWL,N72_PWL,N73_PWL,N74_PWL,N75_PWL,N80_PWL,N85_PWL,N86_PWL,N87_PWL,
            N88_PWL,N89_PWL,N90_PWL,N91_PWL,N96_PWL,N101_PWL,N106_PWL,N111_PWL,N116_PWL,N121_PWL,
            N126_PWL,N130_PWL,N135_PWL,N138_PWL,N143_PWL,N146_PWL,N149_PWL,N152_PWL,N153_PWL,N156_PWL,
            N159_PWL,N165_PWL,N171_PWL,N177_PWL,N183_PWL,N189_PWL,N195_PWL,N201_PWL,N207_PWL,N210_PWL,
            N219_PWL,N228_PWL,N237_PWL,N246_PWL,N255_PWL,N259_PWL,N260_PWL,N261_PWL,N267_PWL,N268_PWL;

      output N388_TERMINATION,N389_TERMINATION,N390_TERMINATION,N391_TERMINATION,N418_TERMINATION,
      N419_TERMINATION,N420_TERMINATION,N421_TERMINATION,N422_TERMINATION,N423_TERMINATION,
      N446_TERMINATION,N447_TERMINATION,N448_TERMINATION,N449_TERMINATION,N450_TERMINATION,
      N767_TERMINATION,N768_TERMINATION,N850_TERMINATION,N863_TERMINATION,N864_TERMINATION,
      N865_TERMINATION,N866_TERMINATION,N874_TERMINATION,N878_TERMINATION,N879_TERMINATION,
      N880_TERMINATION;

      wire GND = 1'b0;
      wire XNOR_1_1_N1_PULSESHAPING_OUT, XNOR_1_2_N1_PULSESHAPING_OUT, XNOR_1_3_N1_PULSESHAPING_OUT, XNOR_1_4_N1_PULSESHAPING_OUT, XNOR_1_5_N1_PULSESHAPING_OUT, XNOR_1_6_N1_PULSESHAPING_OUT;
      NOR2_X1 XNOR_1_1_N1_PULSESHAPING (.ZN (XNOR_1_1_N1_PULSESHAPING_OUT), .A1 (N1_PWL), .A2 (GND));
      NOR2_X1 XNOR_1_2_N1_PULSESHAPING (.ZN (XNOR_1_2_N1_PULSESHAPING_OUT), .A1 (XNOR_1_1_N1_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_3_N1_PULSESHAPING (.ZN (XNOR_1_3_N1_PULSESHAPING_OUT), .A1 (XNOR_1_2_N1_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_4_N1_PULSESHAPING (.ZN (XNOR_1_4_N1_PULSESHAPING_OUT), .A1 (XNOR_1_3_N1_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_5_N1_PULSESHAPING (.ZN (XNOR_1_5_N1_PULSESHAPING_OUT), .A1 (XNOR_1_4_N1_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_6_N1_PULSESHAPING (.ZN (XNOR_1_6_N1_PULSESHAPING_OUT), .A1 (XNOR_1_5_N1_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_7_N1_PULSESHAPING (.ZN (N1), .A1 (XNOR_1_6_N1_PULSESHAPING_OUT), .A2 (GND));

      wire XNOR_1_1_N8_PULSESHAPING_OUT, XNOR_1_2_N8_PULSESHAPING_OUT, XNOR_1_3_N8_PULSESHAPING_OUT, XNOR_1_4_N8_PULSESHAPING_OUT, XNOR_1_5_N8_PULSESHAPING_OUT, XNOR_1_6_N8_PULSESHAPING_OUT;
      NOR2_X1 XNOR_1_1_N8_PULSESHAPING (.ZN (XNOR_1_1_N8_PULSESHAPING_OUT), .A1 (N8_PWL), .A2 (GND));
      NOR2_X1 XNOR_1_2_N8_PULSESHAPING (.ZN (XNOR_1_2_N8_PULSESHAPING_OUT), .A1 (XNOR_1_1_N8_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_3_N8_PULSESHAPING (.ZN (XNOR_1_3_N8_PULSESHAPING_OUT), .A1 (XNOR_1_2_N8_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_4_N8_PULSESHAPING (.ZN (XNOR_1_4_N8_PULSESHAPING_OUT), .A1 (XNOR_1_3_N8_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_5_N8_PULSESHAPING (.ZN (XNOR_1_5_N8_PULSESHAPING_OUT), .A1 (XNOR_1_4_N8_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_6_N8_PULSESHAPING (.ZN (XNOR_1_6_N8_PULSESHAPING_OUT), .A1 (XNOR_1_5_N8_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_7_N8_PULSESHAPING (.ZN (N8), .A1 (XNOR_1_6_N8_PULSESHAPING_OUT), .A2 (GND));

      wire XNOR_1_1_N13_PULSESHAPING_OUT, XNOR_1_2_N13_PULSESHAPING_OUT, XNOR_1_3_N13_PULSESHAPING_OUT, XNOR_1_4_N13_PULSESHAPING_OUT, XNOR_1_5_N13_PULSESHAPING_OUT, XNOR_1_6_N13_PULSESHAPING_OUT;
      NOR2_X1 XNOR_1_1_N13_PULSESHAPING (.ZN (XNOR_1_1_N13_PULSESHAPING_OUT), .A1 (N13_PWL), .A2 (GND));
      NOR2_X1 XNOR_1_2_N13_PULSESHAPING (.ZN (XNOR_1_2_N13_PULSESHAPING_OUT), .A1 (XNOR_1_1_N13_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_3_N13_PULSESHAPING (.ZN (XNOR_1_3_N13_PULSESHAPING_OUT), .A1 (XNOR_1_2_N13_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_4_N13_PULSESHAPING (.ZN (XNOR_1_4_N13_PULSESHAPING_OUT), .A1 (XNOR_1_3_N13_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_5_N13_PULSESHAPING (.ZN (XNOR_1_5_N13_PULSESHAPING_OUT), .A1 (XNOR_1_4_N13_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_6_N13_PULSESHAPING (.ZN (XNOR_1_6_N13_PULSESHAPING_OUT), .A1 (XNOR_1_5_N13_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_7_N13_PULSESHAPING (.ZN (N13), .A1 (XNOR_1_6_N13_PULSESHAPING_OUT), .A2 (GND));

      wire XNOR_1_1_N17_PULSESHAPING_OUT, XNOR_1_2_N17_PULSESHAPING_OUT, XNOR_1_3_N17_PULSESHAPING_OUT, XNOR_1_4_N17_PULSESHAPING_OUT, XNOR_1_5_N17_PULSESHAPING_OUT, XNOR_1_6_N17_PULSESHAPING_OUT;
      NOR2_X1 XNOR_1_1_N17_PULSESHAPING (.ZN (XNOR_1_1_N17_PULSESHAPING_OUT), .A1 (N17_PWL), .A2 (GND));
      NOR2_X1 XNOR_1_2_N17_PULSESHAPING (.ZN (XNOR_1_2_N17_PULSESHAPING_OUT), .A1 (XNOR_1_1_N17_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_3_N17_PULSESHAPING (.ZN (XNOR_1_3_N17_PULSESHAPING_OUT), .A1 (XNOR_1_2_N17_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_4_N17_PULSESHAPING (.ZN (XNOR_1_4_N17_PULSESHAPING_OUT), .A1 (XNOR_1_3_N17_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_5_N17_PULSESHAPING (.ZN (XNOR_1_5_N17_PULSESHAPING_OUT), .A1 (XNOR_1_4_N17_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_6_N17_PULSESHAPING (.ZN (XNOR_1_6_N17_PULSESHAPING_OUT), .A1 (XNOR_1_5_N17_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_7_N17_PULSESHAPING (.ZN (N17), .A1 (XNOR_1_6_N17_PULSESHAPING_OUT), .A2 (GND));

      wire XNOR_1_1_N26_PULSESHAPING_OUT, XNOR_1_2_N26_PULSESHAPING_OUT, XNOR_1_3_N26_PULSESHAPING_OUT, XNOR_1_4_N26_PULSESHAPING_OUT, XNOR_1_5_N26_PULSESHAPING_OUT, XNOR_1_6_N26_PULSESHAPING_OUT;
      NOR2_X1 XNOR_1_1_N26_PULSESHAPING (.ZN (XNOR_1_1_N26_PULSESHAPING_OUT), .A1 (N26_PWL), .A2 (GND));
      NOR2_X1 XNOR_1_2_N26_PULSESHAPING (.ZN (XNOR_1_2_N26_PULSESHAPING_OUT), .A1 (XNOR_1_1_N26_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_3_N26_PULSESHAPING (.ZN (XNOR_1_3_N26_PULSESHAPING_OUT), .A1 (XNOR_1_2_N26_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_4_N26_PULSESHAPING (.ZN (XNOR_1_4_N26_PULSESHAPING_OUT), .A1 (XNOR_1_3_N26_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_5_N26_PULSESHAPING (.ZN (XNOR_1_5_N26_PULSESHAPING_OUT), .A1 (XNOR_1_4_N26_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_6_N26_PULSESHAPING (.ZN (XNOR_1_6_N26_PULSESHAPING_OUT), .A1 (XNOR_1_5_N26_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_7_N26_PULSESHAPING (.ZN (N26), .A1 (XNOR_1_6_N26_PULSESHAPING_OUT), .A2 (GND));

      wire XNOR_1_1_N29_PULSESHAPING_OUT, XNOR_1_2_N29_PULSESHAPING_OUT, XNOR_1_3_N29_PULSESHAPING_OUT, XNOR_1_4_N29_PULSESHAPING_OUT, XNOR_1_5_N29_PULSESHAPING_OUT, XNOR_1_6_N29_PULSESHAPING_OUT;
      NOR2_X1 XNOR_1_1_N29_PULSESHAPING (.ZN (XNOR_1_1_N29_PULSESHAPING_OUT), .A1 (N29_PWL), .A2 (GND));
      NOR2_X1 XNOR_1_2_N29_PULSESHAPING (.ZN (XNOR_1_2_N29_PULSESHAPING_OUT), .A1 (XNOR_1_1_N29_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_3_N29_PULSESHAPING (.ZN (XNOR_1_3_N29_PULSESHAPING_OUT), .A1 (XNOR_1_2_N29_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_4_N29_PULSESHAPING (.ZN (XNOR_1_4_N29_PULSESHAPING_OUT), .A1 (XNOR_1_3_N29_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_5_N29_PULSESHAPING (.ZN (XNOR_1_5_N29_PULSESHAPING_OUT), .A1 (XNOR_1_4_N29_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_6_N29_PULSESHAPING (.ZN (XNOR_1_6_N29_PULSESHAPING_OUT), .A1 (XNOR_1_5_N29_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_7_N29_PULSESHAPING (.ZN (N29), .A1 (XNOR_1_6_N29_PULSESHAPING_OUT), .A2 (GND));

      wire XNOR_1_1_N36_PULSESHAPING_OUT, XNOR_1_2_N36_PULSESHAPING_OUT, XNOR_1_3_N36_PULSESHAPING_OUT, XNOR_1_4_N36_PULSESHAPING_OUT, XNOR_1_5_N36_PULSESHAPING_OUT, XNOR_1_6_N36_PULSESHAPING_OUT;
      NOR2_X1 XNOR_1_1_N36_PULSESHAPING (.ZN (XNOR_1_1_N36_PULSESHAPING_OUT), .A1 (N36_PWL), .A2 (GND));
      NOR2_X1 XNOR_1_2_N36_PULSESHAPING (.ZN (XNOR_1_2_N36_PULSESHAPING_OUT), .A1 (XNOR_1_1_N36_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_3_N36_PULSESHAPING (.ZN (XNOR_1_3_N36_PULSESHAPING_OUT), .A1 (XNOR_1_2_N36_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_4_N36_PULSESHAPING (.ZN (XNOR_1_4_N36_PULSESHAPING_OUT), .A1 (XNOR_1_3_N36_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_5_N36_PULSESHAPING (.ZN (XNOR_1_5_N36_PULSESHAPING_OUT), .A1 (XNOR_1_4_N36_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_6_N36_PULSESHAPING (.ZN (XNOR_1_6_N36_PULSESHAPING_OUT), .A1 (XNOR_1_5_N36_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_7_N36_PULSESHAPING (.ZN (N36), .A1 (XNOR_1_6_N36_PULSESHAPING_OUT), .A2 (GND));

      wire XNOR_1_1_N42_PULSESHAPING_OUT, XNOR_1_2_N42_PULSESHAPING_OUT, XNOR_1_3_N42_PULSESHAPING_OUT, XNOR_1_4_N42_PULSESHAPING_OUT, XNOR_1_5_N42_PULSESHAPING_OUT, XNOR_1_6_N42_PULSESHAPING_OUT;
      NOR2_X1 XNOR_1_1_N42_PULSESHAPING (.ZN (XNOR_1_1_N42_PULSESHAPING_OUT), .A1 (N42_PWL), .A2 (GND));
      NOR2_X1 XNOR_1_2_N42_PULSESHAPING (.ZN (XNOR_1_2_N42_PULSESHAPING_OUT), .A1 (XNOR_1_1_N42_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_3_N42_PULSESHAPING (.ZN (XNOR_1_3_N42_PULSESHAPING_OUT), .A1 (XNOR_1_2_N42_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_4_N42_PULSESHAPING (.ZN (XNOR_1_4_N42_PULSESHAPING_OUT), .A1 (XNOR_1_3_N42_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_5_N42_PULSESHAPING (.ZN (XNOR_1_5_N42_PULSESHAPING_OUT), .A1 (XNOR_1_4_N42_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_6_N42_PULSESHAPING (.ZN (XNOR_1_6_N42_PULSESHAPING_OUT), .A1 (XNOR_1_5_N42_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_7_N42_PULSESHAPING (.ZN (N42), .A1 (XNOR_1_6_N42_PULSESHAPING_OUT), .A2 (GND));

      wire XNOR_1_1_N51_PULSESHAPING_OUT, XNOR_1_2_N51_PULSESHAPING_OUT, XNOR_1_3_N51_PULSESHAPING_OUT, XNOR_1_4_N51_PULSESHAPING_OUT, XNOR_1_5_N51_PULSESHAPING_OUT, XNOR_1_6_N51_PULSESHAPING_OUT;
      NOR2_X1 XNOR_1_1_N51_PULSESHAPING (.ZN (XNOR_1_1_N51_PULSESHAPING_OUT), .A1 (N51_PWL), .A2 (GND));
      NOR2_X1 XNOR_1_2_N51_PULSESHAPING (.ZN (XNOR_1_2_N51_PULSESHAPING_OUT), .A1 (XNOR_1_1_N51_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_3_N51_PULSESHAPING (.ZN (XNOR_1_3_N51_PULSESHAPING_OUT), .A1 (XNOR_1_2_N51_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_4_N51_PULSESHAPING (.ZN (XNOR_1_4_N51_PULSESHAPING_OUT), .A1 (XNOR_1_3_N51_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_5_N51_PULSESHAPING (.ZN (XNOR_1_5_N51_PULSESHAPING_OUT), .A1 (XNOR_1_4_N51_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_6_N51_PULSESHAPING (.ZN (XNOR_1_6_N51_PULSESHAPING_OUT), .A1 (XNOR_1_5_N51_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_7_N51_PULSESHAPING (.ZN (N51), .A1 (XNOR_1_6_N51_PULSESHAPING_OUT), .A2 (GND));

      wire XNOR_1_1_N55_PULSESHAPING_OUT, XNOR_1_2_N55_PULSESHAPING_OUT, XNOR_1_3_N55_PULSESHAPING_OUT, XNOR_1_4_N55_PULSESHAPING_OUT, XNOR_1_5_N55_PULSESHAPING_OUT, XNOR_1_6_N55_PULSESHAPING_OUT;
      NOR2_X1 XNOR_1_1_N55_PULSESHAPING (.ZN (XNOR_1_1_N55_PULSESHAPING_OUT), .A1 (N55_PWL), .A2 (GND));
      NOR2_X1 XNOR_1_2_N55_PULSESHAPING (.ZN (XNOR_1_2_N55_PULSESHAPING_OUT), .A1 (XNOR_1_1_N55_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_3_N55_PULSESHAPING (.ZN (XNOR_1_3_N55_PULSESHAPING_OUT), .A1 (XNOR_1_2_N55_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_4_N55_PULSESHAPING (.ZN (XNOR_1_4_N55_PULSESHAPING_OUT), .A1 (XNOR_1_3_N55_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_5_N55_PULSESHAPING (.ZN (XNOR_1_5_N55_PULSESHAPING_OUT), .A1 (XNOR_1_4_N55_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_6_N55_PULSESHAPING (.ZN (XNOR_1_6_N55_PULSESHAPING_OUT), .A1 (XNOR_1_5_N55_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_7_N55_PULSESHAPING (.ZN (N55), .A1 (XNOR_1_6_N55_PULSESHAPING_OUT), .A2 (GND));

      wire XNOR_1_1_N59_PULSESHAPING_OUT, XNOR_1_2_N59_PULSESHAPING_OUT, XNOR_1_3_N59_PULSESHAPING_OUT, XNOR_1_4_N59_PULSESHAPING_OUT, XNOR_1_5_N59_PULSESHAPING_OUT, XNOR_1_6_N59_PULSESHAPING_OUT;
      NOR2_X1 XNOR_1_1_N59_PULSESHAPING (.ZN (XNOR_1_1_N59_PULSESHAPING_OUT), .A1 (N59_PWL), .A2 (GND));
      NOR2_X1 XNOR_1_2_N59_PULSESHAPING (.ZN (XNOR_1_2_N59_PULSESHAPING_OUT), .A1 (XNOR_1_1_N59_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_3_N59_PULSESHAPING (.ZN (XNOR_1_3_N59_PULSESHAPING_OUT), .A1 (XNOR_1_2_N59_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_4_N59_PULSESHAPING (.ZN (XNOR_1_4_N59_PULSESHAPING_OUT), .A1 (XNOR_1_3_N59_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_5_N59_PULSESHAPING (.ZN (XNOR_1_5_N59_PULSESHAPING_OUT), .A1 (XNOR_1_4_N59_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_6_N59_PULSESHAPING (.ZN (XNOR_1_6_N59_PULSESHAPING_OUT), .A1 (XNOR_1_5_N59_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_7_N59_PULSESHAPING (.ZN (N59), .A1 (XNOR_1_6_N59_PULSESHAPING_OUT), .A2 (GND));

      wire XNOR_1_1_N68_PULSESHAPING_OUT, XNOR_1_2_N68_PULSESHAPING_OUT, XNOR_1_3_N68_PULSESHAPING_OUT, XNOR_1_4_N68_PULSESHAPING_OUT, XNOR_1_5_N68_PULSESHAPING_OUT, XNOR_1_6_N68_PULSESHAPING_OUT;
      NOR2_X1 XNOR_1_1_N68_PULSESHAPING (.ZN (XNOR_1_1_N68_PULSESHAPING_OUT), .A1 (N68_PWL), .A2 (GND));
      NOR2_X1 XNOR_1_2_N68_PULSESHAPING (.ZN (XNOR_1_2_N68_PULSESHAPING_OUT), .A1 (XNOR_1_1_N68_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_3_N68_PULSESHAPING (.ZN (XNOR_1_3_N68_PULSESHAPING_OUT), .A1 (XNOR_1_2_N68_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_4_N68_PULSESHAPING (.ZN (XNOR_1_4_N68_PULSESHAPING_OUT), .A1 (XNOR_1_3_N68_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_5_N68_PULSESHAPING (.ZN (XNOR_1_5_N68_PULSESHAPING_OUT), .A1 (XNOR_1_4_N68_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_6_N68_PULSESHAPING (.ZN (XNOR_1_6_N68_PULSESHAPING_OUT), .A1 (XNOR_1_5_N68_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_7_N68_PULSESHAPING (.ZN (N68), .A1 (XNOR_1_6_N68_PULSESHAPING_OUT), .A2 (GND));

      wire XNOR_1_1_N72_PULSESHAPING_OUT, XNOR_1_2_N72_PULSESHAPING_OUT, XNOR_1_3_N72_PULSESHAPING_OUT, XNOR_1_4_N72_PULSESHAPING_OUT, XNOR_1_5_N72_PULSESHAPING_OUT, XNOR_1_6_N72_PULSESHAPING_OUT;
      NOR2_X1 XNOR_1_1_N72_PULSESHAPING (.ZN (XNOR_1_1_N72_PULSESHAPING_OUT), .A1 (N72_PWL), .A2 (GND));
      NOR2_X1 XNOR_1_2_N72_PULSESHAPING (.ZN (XNOR_1_2_N72_PULSESHAPING_OUT), .A1 (XNOR_1_1_N72_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_3_N72_PULSESHAPING (.ZN (XNOR_1_3_N72_PULSESHAPING_OUT), .A1 (XNOR_1_2_N72_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_4_N72_PULSESHAPING (.ZN (XNOR_1_4_N72_PULSESHAPING_OUT), .A1 (XNOR_1_3_N72_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_5_N72_PULSESHAPING (.ZN (XNOR_1_5_N72_PULSESHAPING_OUT), .A1 (XNOR_1_4_N72_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_6_N72_PULSESHAPING (.ZN (XNOR_1_6_N72_PULSESHAPING_OUT), .A1 (XNOR_1_5_N72_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_7_N72_PULSESHAPING (.ZN (N72), .A1 (XNOR_1_6_N72_PULSESHAPING_OUT), .A2 (GND));

      wire XNOR_1_1_N73_PULSESHAPING_OUT, XNOR_1_2_N73_PULSESHAPING_OUT, XNOR_1_3_N73_PULSESHAPING_OUT, XNOR_1_4_N73_PULSESHAPING_OUT, XNOR_1_5_N73_PULSESHAPING_OUT, XNOR_1_6_N73_PULSESHAPING_OUT;
      NOR2_X1 XNOR_1_1_N73_PULSESHAPING (.ZN (XNOR_1_1_N73_PULSESHAPING_OUT), .A1 (N73_PWL), .A2 (GND));
      NOR2_X1 XNOR_1_2_N73_PULSESHAPING (.ZN (XNOR_1_2_N73_PULSESHAPING_OUT), .A1 (XNOR_1_1_N73_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_3_N73_PULSESHAPING (.ZN (XNOR_1_3_N73_PULSESHAPING_OUT), .A1 (XNOR_1_2_N73_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_4_N73_PULSESHAPING (.ZN (XNOR_1_4_N73_PULSESHAPING_OUT), .A1 (XNOR_1_3_N73_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_5_N73_PULSESHAPING (.ZN (XNOR_1_5_N73_PULSESHAPING_OUT), .A1 (XNOR_1_4_N73_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_6_N73_PULSESHAPING (.ZN (XNOR_1_6_N73_PULSESHAPING_OUT), .A1 (XNOR_1_5_N73_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_7_N73_PULSESHAPING (.ZN (N73), .A1 (XNOR_1_6_N73_PULSESHAPING_OUT), .A2 (GND));

      wire XNOR_1_1_N74_PULSESHAPING_OUT, XNOR_1_2_N74_PULSESHAPING_OUT, XNOR_1_3_N74_PULSESHAPING_OUT, XNOR_1_4_N74_PULSESHAPING_OUT, XNOR_1_5_N74_PULSESHAPING_OUT, XNOR_1_6_N74_PULSESHAPING_OUT;
      NOR2_X1 XNOR_1_1_N74_PULSESHAPING (.ZN (XNOR_1_1_N74_PULSESHAPING_OUT), .A1 (N74_PWL), .A2 (GND));
      NOR2_X1 XNOR_1_2_N74_PULSESHAPING (.ZN (XNOR_1_2_N74_PULSESHAPING_OUT), .A1 (XNOR_1_1_N74_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_3_N74_PULSESHAPING (.ZN (XNOR_1_3_N74_PULSESHAPING_OUT), .A1 (XNOR_1_2_N74_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_4_N74_PULSESHAPING (.ZN (XNOR_1_4_N74_PULSESHAPING_OUT), .A1 (XNOR_1_3_N74_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_5_N74_PULSESHAPING (.ZN (XNOR_1_5_N74_PULSESHAPING_OUT), .A1 (XNOR_1_4_N74_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_6_N74_PULSESHAPING (.ZN (XNOR_1_6_N74_PULSESHAPING_OUT), .A1 (XNOR_1_5_N74_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_7_N74_PULSESHAPING (.ZN (N74), .A1 (XNOR_1_6_N74_PULSESHAPING_OUT), .A2 (GND));

      wire XNOR_1_1_N75_PULSESHAPING_OUT, XNOR_1_2_N75_PULSESHAPING_OUT, XNOR_1_3_N75_PULSESHAPING_OUT, XNOR_1_4_N75_PULSESHAPING_OUT, XNOR_1_5_N75_PULSESHAPING_OUT, XNOR_1_6_N75_PULSESHAPING_OUT;
      NOR2_X1 XNOR_1_1_N75_PULSESHAPING (.ZN (XNOR_1_1_N75_PULSESHAPING_OUT), .A1 (N75_PWL), .A2 (GND));
      NOR2_X1 XNOR_1_2_N75_PULSESHAPING (.ZN (XNOR_1_2_N75_PULSESHAPING_OUT), .A1 (XNOR_1_1_N75_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_3_N75_PULSESHAPING (.ZN (XNOR_1_3_N75_PULSESHAPING_OUT), .A1 (XNOR_1_2_N75_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_4_N75_PULSESHAPING (.ZN (XNOR_1_4_N75_PULSESHAPING_OUT), .A1 (XNOR_1_3_N75_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_5_N75_PULSESHAPING (.ZN (XNOR_1_5_N75_PULSESHAPING_OUT), .A1 (XNOR_1_4_N75_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_6_N75_PULSESHAPING (.ZN (XNOR_1_6_N75_PULSESHAPING_OUT), .A1 (XNOR_1_5_N75_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_7_N75_PULSESHAPING (.ZN (N75), .A1 (XNOR_1_6_N75_PULSESHAPING_OUT), .A2 (GND));

      wire XNOR_1_1_N80_PULSESHAPING_OUT, XNOR_1_2_N80_PULSESHAPING_OUT, XNOR_1_3_N80_PULSESHAPING_OUT, XNOR_1_4_N80_PULSESHAPING_OUT, XNOR_1_5_N80_PULSESHAPING_OUT, XNOR_1_6_N80_PULSESHAPING_OUT;
      NOR2_X1 XNOR_1_1_N80_PULSESHAPING (.ZN (XNOR_1_1_N80_PULSESHAPING_OUT), .A1 (N80_PWL), .A2 (GND));
      NOR2_X1 XNOR_1_2_N80_PULSESHAPING (.ZN (XNOR_1_2_N80_PULSESHAPING_OUT), .A1 (XNOR_1_1_N80_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_3_N80_PULSESHAPING (.ZN (XNOR_1_3_N80_PULSESHAPING_OUT), .A1 (XNOR_1_2_N80_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_4_N80_PULSESHAPING (.ZN (XNOR_1_4_N80_PULSESHAPING_OUT), .A1 (XNOR_1_3_N80_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_5_N80_PULSESHAPING (.ZN (XNOR_1_5_N80_PULSESHAPING_OUT), .A1 (XNOR_1_4_N80_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_6_N80_PULSESHAPING (.ZN (XNOR_1_6_N80_PULSESHAPING_OUT), .A1 (XNOR_1_5_N80_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_7_N80_PULSESHAPING (.ZN (N80), .A1 (XNOR_1_6_N80_PULSESHAPING_OUT), .A2 (GND));

      wire XNOR_1_1_N85_PULSESHAPING_OUT, XNOR_1_2_N85_PULSESHAPING_OUT, XNOR_1_3_N85_PULSESHAPING_OUT, XNOR_1_4_N85_PULSESHAPING_OUT, XNOR_1_5_N85_PULSESHAPING_OUT, XNOR_1_6_N85_PULSESHAPING_OUT;
      NOR2_X1 XNOR_1_1_N85_PULSESHAPING (.ZN (XNOR_1_1_N85_PULSESHAPING_OUT), .A1 (N85_PWL), .A2 (GND));
      NOR2_X1 XNOR_1_2_N85_PULSESHAPING (.ZN (XNOR_1_2_N85_PULSESHAPING_OUT), .A1 (XNOR_1_1_N85_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_3_N85_PULSESHAPING (.ZN (XNOR_1_3_N85_PULSESHAPING_OUT), .A1 (XNOR_1_2_N85_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_4_N85_PULSESHAPING (.ZN (XNOR_1_4_N85_PULSESHAPING_OUT), .A1 (XNOR_1_3_N85_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_5_N85_PULSESHAPING (.ZN (XNOR_1_5_N85_PULSESHAPING_OUT), .A1 (XNOR_1_4_N85_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_6_N85_PULSESHAPING (.ZN (XNOR_1_6_N85_PULSESHAPING_OUT), .A1 (XNOR_1_5_N85_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_7_N85_PULSESHAPING (.ZN (N85), .A1 (XNOR_1_6_N85_PULSESHAPING_OUT), .A2 (GND));

      wire XNOR_1_1_N86_PULSESHAPING_OUT, XNOR_1_2_N86_PULSESHAPING_OUT, XNOR_1_3_N86_PULSESHAPING_OUT, XNOR_1_4_N86_PULSESHAPING_OUT, XNOR_1_5_N86_PULSESHAPING_OUT, XNOR_1_6_N86_PULSESHAPING_OUT;
      NOR2_X1 XNOR_1_1_N86_PULSESHAPING (.ZN (XNOR_1_1_N86_PULSESHAPING_OUT), .A1 (N86_PWL), .A2 (GND));
      NOR2_X1 XNOR_1_2_N86_PULSESHAPING (.ZN (XNOR_1_2_N86_PULSESHAPING_OUT), .A1 (XNOR_1_1_N86_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_3_N86_PULSESHAPING (.ZN (XNOR_1_3_N86_PULSESHAPING_OUT), .A1 (XNOR_1_2_N86_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_4_N86_PULSESHAPING (.ZN (XNOR_1_4_N86_PULSESHAPING_OUT), .A1 (XNOR_1_3_N86_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_5_N86_PULSESHAPING (.ZN (XNOR_1_5_N86_PULSESHAPING_OUT), .A1 (XNOR_1_4_N86_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_6_N86_PULSESHAPING (.ZN (XNOR_1_6_N86_PULSESHAPING_OUT), .A1 (XNOR_1_5_N86_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_7_N86_PULSESHAPING (.ZN (N86), .A1 (XNOR_1_6_N86_PULSESHAPING_OUT), .A2 (GND));

      wire XNOR_1_1_N87_PULSESHAPING_OUT, XNOR_1_2_N87_PULSESHAPING_OUT, XNOR_1_3_N87_PULSESHAPING_OUT, XNOR_1_4_N87_PULSESHAPING_OUT, XNOR_1_5_N87_PULSESHAPING_OUT, XNOR_1_6_N87_PULSESHAPING_OUT;
      NOR2_X1 XNOR_1_1_N87_PULSESHAPING (.ZN (XNOR_1_1_N87_PULSESHAPING_OUT), .A1 (N87_PWL), .A2 (GND));
      NOR2_X1 XNOR_1_2_N87_PULSESHAPING (.ZN (XNOR_1_2_N87_PULSESHAPING_OUT), .A1 (XNOR_1_1_N87_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_3_N87_PULSESHAPING (.ZN (XNOR_1_3_N87_PULSESHAPING_OUT), .A1 (XNOR_1_2_N87_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_4_N87_PULSESHAPING (.ZN (XNOR_1_4_N87_PULSESHAPING_OUT), .A1 (XNOR_1_3_N87_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_5_N87_PULSESHAPING (.ZN (XNOR_1_5_N87_PULSESHAPING_OUT), .A1 (XNOR_1_4_N87_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_6_N87_PULSESHAPING (.ZN (XNOR_1_6_N87_PULSESHAPING_OUT), .A1 (XNOR_1_5_N87_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_7_N87_PULSESHAPING (.ZN (N87), .A1 (XNOR_1_6_N87_PULSESHAPING_OUT), .A2 (GND));

      wire XNOR_1_1_N88_PULSESHAPING_OUT, XNOR_1_2_N88_PULSESHAPING_OUT, XNOR_1_3_N88_PULSESHAPING_OUT, XNOR_1_4_N88_PULSESHAPING_OUT, XNOR_1_5_N88_PULSESHAPING_OUT, XNOR_1_6_N88_PULSESHAPING_OUT;
      NOR2_X1 XNOR_1_1_N88_PULSESHAPING (.ZN (XNOR_1_1_N88_PULSESHAPING_OUT), .A1 (N88_PWL), .A2 (GND));
      NOR2_X1 XNOR_1_2_N88_PULSESHAPING (.ZN (XNOR_1_2_N88_PULSESHAPING_OUT), .A1 (XNOR_1_1_N88_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_3_N88_PULSESHAPING (.ZN (XNOR_1_3_N88_PULSESHAPING_OUT), .A1 (XNOR_1_2_N88_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_4_N88_PULSESHAPING (.ZN (XNOR_1_4_N88_PULSESHAPING_OUT), .A1 (XNOR_1_3_N88_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_5_N88_PULSESHAPING (.ZN (XNOR_1_5_N88_PULSESHAPING_OUT), .A1 (XNOR_1_4_N88_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_6_N88_PULSESHAPING (.ZN (XNOR_1_6_N88_PULSESHAPING_OUT), .A1 (XNOR_1_5_N88_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_7_N88_PULSESHAPING (.ZN (N88), .A1 (XNOR_1_6_N88_PULSESHAPING_OUT), .A2 (GND));

      wire XNOR_1_1_N89_PULSESHAPING_OUT, XNOR_1_2_N89_PULSESHAPING_OUT, XNOR_1_3_N89_PULSESHAPING_OUT, XNOR_1_4_N89_PULSESHAPING_OUT, XNOR_1_5_N89_PULSESHAPING_OUT, XNOR_1_6_N89_PULSESHAPING_OUT;
      NOR2_X1 XNOR_1_1_N89_PULSESHAPING (.ZN (XNOR_1_1_N89_PULSESHAPING_OUT), .A1 (N89_PWL), .A2 (GND));
      NOR2_X1 XNOR_1_2_N89_PULSESHAPING (.ZN (XNOR_1_2_N89_PULSESHAPING_OUT), .A1 (XNOR_1_1_N89_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_3_N89_PULSESHAPING (.ZN (XNOR_1_3_N89_PULSESHAPING_OUT), .A1 (XNOR_1_2_N89_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_4_N89_PULSESHAPING (.ZN (XNOR_1_4_N89_PULSESHAPING_OUT), .A1 (XNOR_1_3_N89_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_5_N89_PULSESHAPING (.ZN (XNOR_1_5_N89_PULSESHAPING_OUT), .A1 (XNOR_1_4_N89_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_6_N89_PULSESHAPING (.ZN (XNOR_1_6_N89_PULSESHAPING_OUT), .A1 (XNOR_1_5_N89_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_7_N89_PULSESHAPING (.ZN (N89), .A1 (XNOR_1_6_N89_PULSESHAPING_OUT), .A2 (GND));

      wire XNOR_1_1_N90_PULSESHAPING_OUT, XNOR_1_2_N90_PULSESHAPING_OUT, XNOR_1_3_N90_PULSESHAPING_OUT, XNOR_1_4_N90_PULSESHAPING_OUT, XNOR_1_5_N90_PULSESHAPING_OUT, XNOR_1_6_N90_PULSESHAPING_OUT;
      NOR2_X1 XNOR_1_1_N90_PULSESHAPING (.ZN (XNOR_1_1_N90_PULSESHAPING_OUT), .A1 (N90_PWL), .A2 (GND));
      NOR2_X1 XNOR_1_2_N90_PULSESHAPING (.ZN (XNOR_1_2_N90_PULSESHAPING_OUT), .A1 (XNOR_1_1_N90_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_3_N90_PULSESHAPING (.ZN (XNOR_1_3_N90_PULSESHAPING_OUT), .A1 (XNOR_1_2_N90_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_4_N90_PULSESHAPING (.ZN (XNOR_1_4_N90_PULSESHAPING_OUT), .A1 (XNOR_1_3_N90_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_5_N90_PULSESHAPING (.ZN (XNOR_1_5_N90_PULSESHAPING_OUT), .A1 (XNOR_1_4_N90_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_6_N90_PULSESHAPING (.ZN (XNOR_1_6_N90_PULSESHAPING_OUT), .A1 (XNOR_1_5_N90_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_7_N90_PULSESHAPING (.ZN (N90), .A1 (XNOR_1_6_N90_PULSESHAPING_OUT), .A2 (GND));

      wire XNOR_1_1_N91_PULSESHAPING_OUT, XNOR_1_2_N91_PULSESHAPING_OUT, XNOR_1_3_N91_PULSESHAPING_OUT, XNOR_1_4_N91_PULSESHAPING_OUT, XNOR_1_5_N91_PULSESHAPING_OUT, XNOR_1_6_N91_PULSESHAPING_OUT;
      NOR2_X1 XNOR_1_1_N91_PULSESHAPING (.ZN (XNOR_1_1_N91_PULSESHAPING_OUT), .A1 (N91_PWL), .A2 (GND));
      NOR2_X1 XNOR_1_2_N91_PULSESHAPING (.ZN (XNOR_1_2_N91_PULSESHAPING_OUT), .A1 (XNOR_1_1_N91_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_3_N91_PULSESHAPING (.ZN (XNOR_1_3_N91_PULSESHAPING_OUT), .A1 (XNOR_1_2_N91_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_4_N91_PULSESHAPING (.ZN (XNOR_1_4_N91_PULSESHAPING_OUT), .A1 (XNOR_1_3_N91_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_5_N91_PULSESHAPING (.ZN (XNOR_1_5_N91_PULSESHAPING_OUT), .A1 (XNOR_1_4_N91_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_6_N91_PULSESHAPING (.ZN (XNOR_1_6_N91_PULSESHAPING_OUT), .A1 (XNOR_1_5_N91_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_7_N91_PULSESHAPING (.ZN (N91), .A1 (XNOR_1_6_N91_PULSESHAPING_OUT), .A2 (GND));

      wire XNOR_1_1_N96_PULSESHAPING_OUT, XNOR_1_2_N96_PULSESHAPING_OUT, XNOR_1_3_N96_PULSESHAPING_OUT, XNOR_1_4_N96_PULSESHAPING_OUT, XNOR_1_5_N96_PULSESHAPING_OUT, XNOR_1_6_N96_PULSESHAPING_OUT;
      NOR2_X1 XNOR_1_1_N96_PULSESHAPING (.ZN (XNOR_1_1_N96_PULSESHAPING_OUT), .A1 (N96_PWL), .A2 (GND));
      NOR2_X1 XNOR_1_2_N96_PULSESHAPING (.ZN (XNOR_1_2_N96_PULSESHAPING_OUT), .A1 (XNOR_1_1_N96_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_3_N96_PULSESHAPING (.ZN (XNOR_1_3_N96_PULSESHAPING_OUT), .A1 (XNOR_1_2_N96_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_4_N96_PULSESHAPING (.ZN (XNOR_1_4_N96_PULSESHAPING_OUT), .A1 (XNOR_1_3_N96_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_5_N96_PULSESHAPING (.ZN (XNOR_1_5_N96_PULSESHAPING_OUT), .A1 (XNOR_1_4_N96_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_6_N96_PULSESHAPING (.ZN (XNOR_1_6_N96_PULSESHAPING_OUT), .A1 (XNOR_1_5_N96_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_7_N96_PULSESHAPING (.ZN (N96), .A1 (XNOR_1_6_N96_PULSESHAPING_OUT), .A2 (GND));

      wire XNOR_1_1_N101_PULSESHAPING_OUT, XNOR_1_2_N101_PULSESHAPING_OUT, XNOR_1_3_N101_PULSESHAPING_OUT, XNOR_1_4_N101_PULSESHAPING_OUT, XNOR_1_5_N101_PULSESHAPING_OUT, XNOR_1_6_N101_PULSESHAPING_OUT;
      NOR2_X1 XNOR_1_1_N101_PULSESHAPING (.ZN (XNOR_1_1_N101_PULSESHAPING_OUT), .A1 (N101_PWL), .A2 (GND));
      NOR2_X1 XNOR_1_2_N101_PULSESHAPING (.ZN (XNOR_1_2_N101_PULSESHAPING_OUT), .A1 (XNOR_1_1_N101_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_3_N101_PULSESHAPING (.ZN (XNOR_1_3_N101_PULSESHAPING_OUT), .A1 (XNOR_1_2_N101_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_4_N101_PULSESHAPING (.ZN (XNOR_1_4_N101_PULSESHAPING_OUT), .A1 (XNOR_1_3_N101_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_5_N101_PULSESHAPING (.ZN (XNOR_1_5_N101_PULSESHAPING_OUT), .A1 (XNOR_1_4_N101_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_6_N101_PULSESHAPING (.ZN (XNOR_1_6_N101_PULSESHAPING_OUT), .A1 (XNOR_1_5_N101_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_7_N101_PULSESHAPING (.ZN (N101), .A1 (XNOR_1_6_N101_PULSESHAPING_OUT), .A2 (GND));

      wire XNOR_1_1_N106_PULSESHAPING_OUT, XNOR_1_2_N106_PULSESHAPING_OUT, XNOR_1_3_N106_PULSESHAPING_OUT, XNOR_1_4_N106_PULSESHAPING_OUT, XNOR_1_5_N106_PULSESHAPING_OUT, XNOR_1_6_N106_PULSESHAPING_OUT;
      NOR2_X1 XNOR_1_1_N106_PULSESHAPING (.ZN (XNOR_1_1_N106_PULSESHAPING_OUT), .A1 (N106_PWL), .A2 (GND));
      NOR2_X1 XNOR_1_2_N106_PULSESHAPING (.ZN (XNOR_1_2_N106_PULSESHAPING_OUT), .A1 (XNOR_1_1_N106_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_3_N106_PULSESHAPING (.ZN (XNOR_1_3_N106_PULSESHAPING_OUT), .A1 (XNOR_1_2_N106_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_4_N106_PULSESHAPING (.ZN (XNOR_1_4_N106_PULSESHAPING_OUT), .A1 (XNOR_1_3_N106_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_5_N106_PULSESHAPING (.ZN (XNOR_1_5_N106_PULSESHAPING_OUT), .A1 (XNOR_1_4_N106_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_6_N106_PULSESHAPING (.ZN (XNOR_1_6_N106_PULSESHAPING_OUT), .A1 (XNOR_1_5_N106_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_7_N106_PULSESHAPING (.ZN (N106), .A1 (XNOR_1_6_N106_PULSESHAPING_OUT), .A2 (GND));

      wire XNOR_1_1_N111_PULSESHAPING_OUT, XNOR_1_2_N111_PULSESHAPING_OUT, XNOR_1_3_N111_PULSESHAPING_OUT, XNOR_1_4_N111_PULSESHAPING_OUT, XNOR_1_5_N111_PULSESHAPING_OUT, XNOR_1_6_N111_PULSESHAPING_OUT;
      NOR2_X1 XNOR_1_1_N111_PULSESHAPING (.ZN (XNOR_1_1_N111_PULSESHAPING_OUT), .A1 (N111_PWL), .A2 (GND));
      NOR2_X1 XNOR_1_2_N111_PULSESHAPING (.ZN (XNOR_1_2_N111_PULSESHAPING_OUT), .A1 (XNOR_1_1_N111_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_3_N111_PULSESHAPING (.ZN (XNOR_1_3_N111_PULSESHAPING_OUT), .A1 (XNOR_1_2_N111_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_4_N111_PULSESHAPING (.ZN (XNOR_1_4_N111_PULSESHAPING_OUT), .A1 (XNOR_1_3_N111_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_5_N111_PULSESHAPING (.ZN (XNOR_1_5_N111_PULSESHAPING_OUT), .A1 (XNOR_1_4_N111_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_6_N111_PULSESHAPING (.ZN (XNOR_1_6_N111_PULSESHAPING_OUT), .A1 (XNOR_1_5_N111_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_7_N111_PULSESHAPING (.ZN (N111), .A1 (XNOR_1_6_N111_PULSESHAPING_OUT), .A2 (GND));

      wire XNOR_1_1_N116_PULSESHAPING_OUT, XNOR_1_2_N116_PULSESHAPING_OUT, XNOR_1_3_N116_PULSESHAPING_OUT, XNOR_1_4_N116_PULSESHAPING_OUT, XNOR_1_5_N116_PULSESHAPING_OUT, XNOR_1_6_N116_PULSESHAPING_OUT;
      NOR2_X1 XNOR_1_1_N116_PULSESHAPING (.ZN (XNOR_1_1_N116_PULSESHAPING_OUT), .A1 (N116_PWL), .A2 (GND));
      NOR2_X1 XNOR_1_2_N116_PULSESHAPING (.ZN (XNOR_1_2_N116_PULSESHAPING_OUT), .A1 (XNOR_1_1_N116_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_3_N116_PULSESHAPING (.ZN (XNOR_1_3_N116_PULSESHAPING_OUT), .A1 (XNOR_1_2_N116_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_4_N116_PULSESHAPING (.ZN (XNOR_1_4_N116_PULSESHAPING_OUT), .A1 (XNOR_1_3_N116_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_5_N116_PULSESHAPING (.ZN (XNOR_1_5_N116_PULSESHAPING_OUT), .A1 (XNOR_1_4_N116_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_6_N116_PULSESHAPING (.ZN (XNOR_1_6_N116_PULSESHAPING_OUT), .A1 (XNOR_1_5_N116_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_7_N116_PULSESHAPING (.ZN (N116), .A1 (XNOR_1_6_N116_PULSESHAPING_OUT), .A2 (GND));

      wire XNOR_1_1_N121_PULSESHAPING_OUT, XNOR_1_2_N121_PULSESHAPING_OUT, XNOR_1_3_N121_PULSESHAPING_OUT, XNOR_1_4_N121_PULSESHAPING_OUT, XNOR_1_5_N121_PULSESHAPING_OUT, XNOR_1_6_N121_PULSESHAPING_OUT;
      NOR2_X1 XNOR_1_1_N121_PULSESHAPING (.ZN (XNOR_1_1_N121_PULSESHAPING_OUT), .A1 (N121_PWL), .A2 (GND));
      NOR2_X1 XNOR_1_2_N121_PULSESHAPING (.ZN (XNOR_1_2_N121_PULSESHAPING_OUT), .A1 (XNOR_1_1_N121_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_3_N121_PULSESHAPING (.ZN (XNOR_1_3_N121_PULSESHAPING_OUT), .A1 (XNOR_1_2_N121_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_4_N121_PULSESHAPING (.ZN (XNOR_1_4_N121_PULSESHAPING_OUT), .A1 (XNOR_1_3_N121_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_5_N121_PULSESHAPING (.ZN (XNOR_1_5_N121_PULSESHAPING_OUT), .A1 (XNOR_1_4_N121_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_6_N121_PULSESHAPING (.ZN (XNOR_1_6_N121_PULSESHAPING_OUT), .A1 (XNOR_1_5_N121_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_7_N121_PULSESHAPING (.ZN (N121), .A1 (XNOR_1_6_N121_PULSESHAPING_OUT), .A2 (GND));

      wire XNOR_1_1_N126_PULSESHAPING_OUT, XNOR_1_2_N126_PULSESHAPING_OUT, XNOR_1_3_N126_PULSESHAPING_OUT, XNOR_1_4_N126_PULSESHAPING_OUT, XNOR_1_5_N126_PULSESHAPING_OUT, XNOR_1_6_N126_PULSESHAPING_OUT;
      NOR2_X1 XNOR_1_1_N126_PULSESHAPING (.ZN (XNOR_1_1_N126_PULSESHAPING_OUT), .A1 (N126_PWL), .A2 (GND));
      NOR2_X1 XNOR_1_2_N126_PULSESHAPING (.ZN (XNOR_1_2_N126_PULSESHAPING_OUT), .A1 (XNOR_1_1_N126_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_3_N126_PULSESHAPING (.ZN (XNOR_1_3_N126_PULSESHAPING_OUT), .A1 (XNOR_1_2_N126_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_4_N126_PULSESHAPING (.ZN (XNOR_1_4_N126_PULSESHAPING_OUT), .A1 (XNOR_1_3_N126_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_5_N126_PULSESHAPING (.ZN (XNOR_1_5_N126_PULSESHAPING_OUT), .A1 (XNOR_1_4_N126_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_6_N126_PULSESHAPING (.ZN (XNOR_1_6_N126_PULSESHAPING_OUT), .A1 (XNOR_1_5_N126_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_7_N126_PULSESHAPING (.ZN (N126), .A1 (XNOR_1_6_N126_PULSESHAPING_OUT), .A2 (GND));

      wire XNOR_1_1_N130_PULSESHAPING_OUT, XNOR_1_2_N130_PULSESHAPING_OUT, XNOR_1_3_N130_PULSESHAPING_OUT, XNOR_1_4_N130_PULSESHAPING_OUT, XNOR_1_5_N130_PULSESHAPING_OUT, XNOR_1_6_N130_PULSESHAPING_OUT;
      NOR2_X1 XNOR_1_1_N130_PULSESHAPING (.ZN (XNOR_1_1_N130_PULSESHAPING_OUT), .A1 (N130_PWL), .A2 (GND));
      NOR2_X1 XNOR_1_2_N130_PULSESHAPING (.ZN (XNOR_1_2_N130_PULSESHAPING_OUT), .A1 (XNOR_1_1_N130_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_3_N130_PULSESHAPING (.ZN (XNOR_1_3_N130_PULSESHAPING_OUT), .A1 (XNOR_1_2_N130_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_4_N130_PULSESHAPING (.ZN (XNOR_1_4_N130_PULSESHAPING_OUT), .A1 (XNOR_1_3_N130_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_5_N130_PULSESHAPING (.ZN (XNOR_1_5_N130_PULSESHAPING_OUT), .A1 (XNOR_1_4_N130_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_6_N130_PULSESHAPING (.ZN (XNOR_1_6_N130_PULSESHAPING_OUT), .A1 (XNOR_1_5_N130_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_7_N130_PULSESHAPING (.ZN (N130), .A1 (XNOR_1_6_N130_PULSESHAPING_OUT), .A2 (GND));

      wire XNOR_1_1_N135_PULSESHAPING_OUT, XNOR_1_2_N135_PULSESHAPING_OUT, XNOR_1_3_N135_PULSESHAPING_OUT, XNOR_1_4_N135_PULSESHAPING_OUT, XNOR_1_5_N135_PULSESHAPING_OUT, XNOR_1_6_N135_PULSESHAPING_OUT;
      NOR2_X1 XNOR_1_1_N135_PULSESHAPING (.ZN (XNOR_1_1_N135_PULSESHAPING_OUT), .A1 (N135_PWL), .A2 (GND));
      NOR2_X1 XNOR_1_2_N135_PULSESHAPING (.ZN (XNOR_1_2_N135_PULSESHAPING_OUT), .A1 (XNOR_1_1_N135_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_3_N135_PULSESHAPING (.ZN (XNOR_1_3_N135_PULSESHAPING_OUT), .A1 (XNOR_1_2_N135_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_4_N135_PULSESHAPING (.ZN (XNOR_1_4_N135_PULSESHAPING_OUT), .A1 (XNOR_1_3_N135_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_5_N135_PULSESHAPING (.ZN (XNOR_1_5_N135_PULSESHAPING_OUT), .A1 (XNOR_1_4_N135_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_6_N135_PULSESHAPING (.ZN (XNOR_1_6_N135_PULSESHAPING_OUT), .A1 (XNOR_1_5_N135_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_7_N135_PULSESHAPING (.ZN (N135), .A1 (XNOR_1_6_N135_PULSESHAPING_OUT), .A2 (GND));

      wire XNOR_1_1_N138_PULSESHAPING_OUT, XNOR_1_2_N138_PULSESHAPING_OUT, XNOR_1_3_N138_PULSESHAPING_OUT, XNOR_1_4_N138_PULSESHAPING_OUT, XNOR_1_5_N138_PULSESHAPING_OUT, XNOR_1_6_N138_PULSESHAPING_OUT;
      NOR2_X1 XNOR_1_1_N138_PULSESHAPING (.ZN (XNOR_1_1_N138_PULSESHAPING_OUT), .A1 (N138_PWL), .A2 (GND));
      NOR2_X1 XNOR_1_2_N138_PULSESHAPING (.ZN (XNOR_1_2_N138_PULSESHAPING_OUT), .A1 (XNOR_1_1_N138_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_3_N138_PULSESHAPING (.ZN (XNOR_1_3_N138_PULSESHAPING_OUT), .A1 (XNOR_1_2_N138_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_4_N138_PULSESHAPING (.ZN (XNOR_1_4_N138_PULSESHAPING_OUT), .A1 (XNOR_1_3_N138_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_5_N138_PULSESHAPING (.ZN (XNOR_1_5_N138_PULSESHAPING_OUT), .A1 (XNOR_1_4_N138_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_6_N138_PULSESHAPING (.ZN (XNOR_1_6_N138_PULSESHAPING_OUT), .A1 (XNOR_1_5_N138_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_7_N138_PULSESHAPING (.ZN (N138), .A1 (XNOR_1_6_N138_PULSESHAPING_OUT), .A2 (GND));

      wire XNOR_1_1_N143_PULSESHAPING_OUT, XNOR_1_2_N143_PULSESHAPING_OUT, XNOR_1_3_N143_PULSESHAPING_OUT, XNOR_1_4_N143_PULSESHAPING_OUT, XNOR_1_5_N143_PULSESHAPING_OUT, XNOR_1_6_N143_PULSESHAPING_OUT;
      NOR2_X1 XNOR_1_1_N143_PULSESHAPING (.ZN (XNOR_1_1_N143_PULSESHAPING_OUT), .A1 (N143_PWL), .A2 (GND));
      NOR2_X1 XNOR_1_2_N143_PULSESHAPING (.ZN (XNOR_1_2_N143_PULSESHAPING_OUT), .A1 (XNOR_1_1_N143_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_3_N143_PULSESHAPING (.ZN (XNOR_1_3_N143_PULSESHAPING_OUT), .A1 (XNOR_1_2_N143_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_4_N143_PULSESHAPING (.ZN (XNOR_1_4_N143_PULSESHAPING_OUT), .A1 (XNOR_1_3_N143_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_5_N143_PULSESHAPING (.ZN (XNOR_1_5_N143_PULSESHAPING_OUT), .A1 (XNOR_1_4_N143_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_6_N143_PULSESHAPING (.ZN (XNOR_1_6_N143_PULSESHAPING_OUT), .A1 (XNOR_1_5_N143_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_7_N143_PULSESHAPING (.ZN (N143), .A1 (XNOR_1_6_N143_PULSESHAPING_OUT), .A2 (GND));

      wire XNOR_1_1_N146_PULSESHAPING_OUT, XNOR_1_2_N146_PULSESHAPING_OUT, XNOR_1_3_N146_PULSESHAPING_OUT, XNOR_1_4_N146_PULSESHAPING_OUT, XNOR_1_5_N146_PULSESHAPING_OUT, XNOR_1_6_N146_PULSESHAPING_OUT;
      NOR2_X1 XNOR_1_1_N146_PULSESHAPING (.ZN (XNOR_1_1_N146_PULSESHAPING_OUT), .A1 (N146_PWL), .A2 (GND));
      NOR2_X1 XNOR_1_2_N146_PULSESHAPING (.ZN (XNOR_1_2_N146_PULSESHAPING_OUT), .A1 (XNOR_1_1_N146_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_3_N146_PULSESHAPING (.ZN (XNOR_1_3_N146_PULSESHAPING_OUT), .A1 (XNOR_1_2_N146_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_4_N146_PULSESHAPING (.ZN (XNOR_1_4_N146_PULSESHAPING_OUT), .A1 (XNOR_1_3_N146_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_5_N146_PULSESHAPING (.ZN (XNOR_1_5_N146_PULSESHAPING_OUT), .A1 (XNOR_1_4_N146_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_6_N146_PULSESHAPING (.ZN (XNOR_1_6_N146_PULSESHAPING_OUT), .A1 (XNOR_1_5_N146_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_7_N146_PULSESHAPING (.ZN (N146), .A1 (XNOR_1_6_N146_PULSESHAPING_OUT), .A2 (GND));

      wire XNOR_1_1_N149_PULSESHAPING_OUT, XNOR_1_2_N149_PULSESHAPING_OUT, XNOR_1_3_N149_PULSESHAPING_OUT, XNOR_1_4_N149_PULSESHAPING_OUT, XNOR_1_5_N149_PULSESHAPING_OUT, XNOR_1_6_N149_PULSESHAPING_OUT;
      NOR2_X1 XNOR_1_1_N149_PULSESHAPING (.ZN (XNOR_1_1_N149_PULSESHAPING_OUT), .A1 (N149_PWL), .A2 (GND));
      NOR2_X1 XNOR_1_2_N149_PULSESHAPING (.ZN (XNOR_1_2_N149_PULSESHAPING_OUT), .A1 (XNOR_1_1_N149_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_3_N149_PULSESHAPING (.ZN (XNOR_1_3_N149_PULSESHAPING_OUT), .A1 (XNOR_1_2_N149_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_4_N149_PULSESHAPING (.ZN (XNOR_1_4_N149_PULSESHAPING_OUT), .A1 (XNOR_1_3_N149_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_5_N149_PULSESHAPING (.ZN (XNOR_1_5_N149_PULSESHAPING_OUT), .A1 (XNOR_1_4_N149_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_6_N149_PULSESHAPING (.ZN (XNOR_1_6_N149_PULSESHAPING_OUT), .A1 (XNOR_1_5_N149_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_7_N149_PULSESHAPING (.ZN (N149), .A1 (XNOR_1_6_N149_PULSESHAPING_OUT), .A2 (GND));

      wire XNOR_1_1_N152_PULSESHAPING_OUT, XNOR_1_2_N152_PULSESHAPING_OUT, XNOR_1_3_N152_PULSESHAPING_OUT, XNOR_1_4_N152_PULSESHAPING_OUT, XNOR_1_5_N152_PULSESHAPING_OUT, XNOR_1_6_N152_PULSESHAPING_OUT;
      NOR2_X1 XNOR_1_1_N152_PULSESHAPING (.ZN (XNOR_1_1_N152_PULSESHAPING_OUT), .A1 (N152_PWL), .A2 (GND));
      NOR2_X1 XNOR_1_2_N152_PULSESHAPING (.ZN (XNOR_1_2_N152_PULSESHAPING_OUT), .A1 (XNOR_1_1_N152_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_3_N152_PULSESHAPING (.ZN (XNOR_1_3_N152_PULSESHAPING_OUT), .A1 (XNOR_1_2_N152_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_4_N152_PULSESHAPING (.ZN (XNOR_1_4_N152_PULSESHAPING_OUT), .A1 (XNOR_1_3_N152_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_5_N152_PULSESHAPING (.ZN (XNOR_1_5_N152_PULSESHAPING_OUT), .A1 (XNOR_1_4_N152_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_6_N152_PULSESHAPING (.ZN (XNOR_1_6_N152_PULSESHAPING_OUT), .A1 (XNOR_1_5_N152_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_7_N152_PULSESHAPING (.ZN (N152), .A1 (XNOR_1_6_N152_PULSESHAPING_OUT), .A2 (GND));

      wire XNOR_1_1_N153_PULSESHAPING_OUT, XNOR_1_2_N153_PULSESHAPING_OUT, XNOR_1_3_N153_PULSESHAPING_OUT, XNOR_1_4_N153_PULSESHAPING_OUT, XNOR_1_5_N153_PULSESHAPING_OUT, XNOR_1_6_N153_PULSESHAPING_OUT;
      NOR2_X1 XNOR_1_1_N153_PULSESHAPING (.ZN (XNOR_1_1_N153_PULSESHAPING_OUT), .A1 (N153_PWL), .A2 (GND));
      NOR2_X1 XNOR_1_2_N153_PULSESHAPING (.ZN (XNOR_1_2_N153_PULSESHAPING_OUT), .A1 (XNOR_1_1_N153_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_3_N153_PULSESHAPING (.ZN (XNOR_1_3_N153_PULSESHAPING_OUT), .A1 (XNOR_1_2_N153_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_4_N153_PULSESHAPING (.ZN (XNOR_1_4_N153_PULSESHAPING_OUT), .A1 (XNOR_1_3_N153_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_5_N153_PULSESHAPING (.ZN (XNOR_1_5_N153_PULSESHAPING_OUT), .A1 (XNOR_1_4_N153_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_6_N153_PULSESHAPING (.ZN (XNOR_1_6_N153_PULSESHAPING_OUT), .A1 (XNOR_1_5_N153_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_7_N153_PULSESHAPING (.ZN (N153), .A1 (XNOR_1_6_N153_PULSESHAPING_OUT), .A2 (GND));

      wire XNOR_1_1_N156_PULSESHAPING_OUT, XNOR_1_2_N156_PULSESHAPING_OUT, XNOR_1_3_N156_PULSESHAPING_OUT, XNOR_1_4_N156_PULSESHAPING_OUT, XNOR_1_5_N156_PULSESHAPING_OUT, XNOR_1_6_N156_PULSESHAPING_OUT;
      NOR2_X1 XNOR_1_1_N156_PULSESHAPING (.ZN (XNOR_1_1_N156_PULSESHAPING_OUT), .A1 (N156_PWL), .A2 (GND));
      NOR2_X1 XNOR_1_2_N156_PULSESHAPING (.ZN (XNOR_1_2_N156_PULSESHAPING_OUT), .A1 (XNOR_1_1_N156_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_3_N156_PULSESHAPING (.ZN (XNOR_1_3_N156_PULSESHAPING_OUT), .A1 (XNOR_1_2_N156_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_4_N156_PULSESHAPING (.ZN (XNOR_1_4_N156_PULSESHAPING_OUT), .A1 (XNOR_1_3_N156_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_5_N156_PULSESHAPING (.ZN (XNOR_1_5_N156_PULSESHAPING_OUT), .A1 (XNOR_1_4_N156_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_6_N156_PULSESHAPING (.ZN (XNOR_1_6_N156_PULSESHAPING_OUT), .A1 (XNOR_1_5_N156_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_7_N156_PULSESHAPING (.ZN (N156), .A1 (XNOR_1_6_N156_PULSESHAPING_OUT), .A2 (GND));

      wire XNOR_1_1_N159_PULSESHAPING_OUT, XNOR_1_2_N159_PULSESHAPING_OUT, XNOR_1_3_N159_PULSESHAPING_OUT, XNOR_1_4_N159_PULSESHAPING_OUT, XNOR_1_5_N159_PULSESHAPING_OUT, XNOR_1_6_N159_PULSESHAPING_OUT;
      NOR2_X1 XNOR_1_1_N159_PULSESHAPING (.ZN (XNOR_1_1_N159_PULSESHAPING_OUT), .A1 (N159_PWL), .A2 (GND));
      NOR2_X1 XNOR_1_2_N159_PULSESHAPING (.ZN (XNOR_1_2_N159_PULSESHAPING_OUT), .A1 (XNOR_1_1_N159_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_3_N159_PULSESHAPING (.ZN (XNOR_1_3_N159_PULSESHAPING_OUT), .A1 (XNOR_1_2_N159_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_4_N159_PULSESHAPING (.ZN (XNOR_1_4_N159_PULSESHAPING_OUT), .A1 (XNOR_1_3_N159_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_5_N159_PULSESHAPING (.ZN (XNOR_1_5_N159_PULSESHAPING_OUT), .A1 (XNOR_1_4_N159_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_6_N159_PULSESHAPING (.ZN (XNOR_1_6_N159_PULSESHAPING_OUT), .A1 (XNOR_1_5_N159_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_7_N159_PULSESHAPING (.ZN (N159), .A1 (XNOR_1_6_N159_PULSESHAPING_OUT), .A2 (GND));

      wire XNOR_1_1_N165_PULSESHAPING_OUT, XNOR_1_2_N165_PULSESHAPING_OUT, XNOR_1_3_N165_PULSESHAPING_OUT, XNOR_1_4_N165_PULSESHAPING_OUT, XNOR_1_5_N165_PULSESHAPING_OUT, XNOR_1_6_N165_PULSESHAPING_OUT;
      NOR2_X1 XNOR_1_1_N165_PULSESHAPING (.ZN (XNOR_1_1_N165_PULSESHAPING_OUT), .A1 (N165_PWL), .A2 (GND));
      NOR2_X1 XNOR_1_2_N165_PULSESHAPING (.ZN (XNOR_1_2_N165_PULSESHAPING_OUT), .A1 (XNOR_1_1_N165_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_3_N165_PULSESHAPING (.ZN (XNOR_1_3_N165_PULSESHAPING_OUT), .A1 (XNOR_1_2_N165_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_4_N165_PULSESHAPING (.ZN (XNOR_1_4_N165_PULSESHAPING_OUT), .A1 (XNOR_1_3_N165_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_5_N165_PULSESHAPING (.ZN (XNOR_1_5_N165_PULSESHAPING_OUT), .A1 (XNOR_1_4_N165_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_6_N165_PULSESHAPING (.ZN (XNOR_1_6_N165_PULSESHAPING_OUT), .A1 (XNOR_1_5_N165_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_7_N165_PULSESHAPING (.ZN (N165), .A1 (XNOR_1_6_N165_PULSESHAPING_OUT), .A2 (GND));

      wire XNOR_1_1_N171_PULSESHAPING_OUT, XNOR_1_2_N171_PULSESHAPING_OUT, XNOR_1_3_N171_PULSESHAPING_OUT, XNOR_1_4_N171_PULSESHAPING_OUT, XNOR_1_5_N171_PULSESHAPING_OUT, XNOR_1_6_N171_PULSESHAPING_OUT;
      NOR2_X1 XNOR_1_1_N171_PULSESHAPING (.ZN (XNOR_1_1_N171_PULSESHAPING_OUT), .A1 (N171_PWL), .A2 (GND));
      NOR2_X1 XNOR_1_2_N171_PULSESHAPING (.ZN (XNOR_1_2_N171_PULSESHAPING_OUT), .A1 (XNOR_1_1_N171_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_3_N171_PULSESHAPING (.ZN (XNOR_1_3_N171_PULSESHAPING_OUT), .A1 (XNOR_1_2_N171_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_4_N171_PULSESHAPING (.ZN (XNOR_1_4_N171_PULSESHAPING_OUT), .A1 (XNOR_1_3_N171_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_5_N171_PULSESHAPING (.ZN (XNOR_1_5_N171_PULSESHAPING_OUT), .A1 (XNOR_1_4_N171_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_6_N171_PULSESHAPING (.ZN (XNOR_1_6_N171_PULSESHAPING_OUT), .A1 (XNOR_1_5_N171_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_7_N171_PULSESHAPING (.ZN (N171), .A1 (XNOR_1_6_N171_PULSESHAPING_OUT), .A2 (GND));

      wire XNOR_1_1_N177_PULSESHAPING_OUT, XNOR_1_2_N177_PULSESHAPING_OUT, XNOR_1_3_N177_PULSESHAPING_OUT, XNOR_1_4_N177_PULSESHAPING_OUT, XNOR_1_5_N177_PULSESHAPING_OUT, XNOR_1_6_N177_PULSESHAPING_OUT;
      NOR2_X1 XNOR_1_1_N177_PULSESHAPING (.ZN (XNOR_1_1_N177_PULSESHAPING_OUT), .A1 (N177_PWL), .A2 (GND));
      NOR2_X1 XNOR_1_2_N177_PULSESHAPING (.ZN (XNOR_1_2_N177_PULSESHAPING_OUT), .A1 (XNOR_1_1_N177_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_3_N177_PULSESHAPING (.ZN (XNOR_1_3_N177_PULSESHAPING_OUT), .A1 (XNOR_1_2_N177_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_4_N177_PULSESHAPING (.ZN (XNOR_1_4_N177_PULSESHAPING_OUT), .A1 (XNOR_1_3_N177_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_5_N177_PULSESHAPING (.ZN (XNOR_1_5_N177_PULSESHAPING_OUT), .A1 (XNOR_1_4_N177_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_6_N177_PULSESHAPING (.ZN (XNOR_1_6_N177_PULSESHAPING_OUT), .A1 (XNOR_1_5_N177_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_7_N177_PULSESHAPING (.ZN (N177), .A1 (XNOR_1_6_N177_PULSESHAPING_OUT), .A2 (GND));

      wire XNOR_1_1_N183_PULSESHAPING_OUT, XNOR_1_2_N183_PULSESHAPING_OUT, XNOR_1_3_N183_PULSESHAPING_OUT, XNOR_1_4_N183_PULSESHAPING_OUT, XNOR_1_5_N183_PULSESHAPING_OUT, XNOR_1_6_N183_PULSESHAPING_OUT;
      NOR2_X1 XNOR_1_1_N183_PULSESHAPING (.ZN (XNOR_1_1_N183_PULSESHAPING_OUT), .A1 (N183_PWL), .A2 (GND));
      NOR2_X1 XNOR_1_2_N183_PULSESHAPING (.ZN (XNOR_1_2_N183_PULSESHAPING_OUT), .A1 (XNOR_1_1_N183_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_3_N183_PULSESHAPING (.ZN (XNOR_1_3_N183_PULSESHAPING_OUT), .A1 (XNOR_1_2_N183_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_4_N183_PULSESHAPING (.ZN (XNOR_1_4_N183_PULSESHAPING_OUT), .A1 (XNOR_1_3_N183_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_5_N183_PULSESHAPING (.ZN (XNOR_1_5_N183_PULSESHAPING_OUT), .A1 (XNOR_1_4_N183_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_6_N183_PULSESHAPING (.ZN (XNOR_1_6_N183_PULSESHAPING_OUT), .A1 (XNOR_1_5_N183_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_7_N183_PULSESHAPING (.ZN (N183), .A1 (XNOR_1_6_N183_PULSESHAPING_OUT), .A2 (GND));

      wire XNOR_1_1_N189_PULSESHAPING_OUT, XNOR_1_2_N189_PULSESHAPING_OUT, XNOR_1_3_N189_PULSESHAPING_OUT, XNOR_1_4_N189_PULSESHAPING_OUT, XNOR_1_5_N189_PULSESHAPING_OUT, XNOR_1_6_N189_PULSESHAPING_OUT;
      NOR2_X1 XNOR_1_1_N189_PULSESHAPING (.ZN (XNOR_1_1_N189_PULSESHAPING_OUT), .A1 (N189_PWL), .A2 (GND));
      NOR2_X1 XNOR_1_2_N189_PULSESHAPING (.ZN (XNOR_1_2_N189_PULSESHAPING_OUT), .A1 (XNOR_1_1_N189_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_3_N189_PULSESHAPING (.ZN (XNOR_1_3_N189_PULSESHAPING_OUT), .A1 (XNOR_1_2_N189_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_4_N189_PULSESHAPING (.ZN (XNOR_1_4_N189_PULSESHAPING_OUT), .A1 (XNOR_1_3_N189_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_5_N189_PULSESHAPING (.ZN (XNOR_1_5_N189_PULSESHAPING_OUT), .A1 (XNOR_1_4_N189_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_6_N189_PULSESHAPING (.ZN (XNOR_1_6_N189_PULSESHAPING_OUT), .A1 (XNOR_1_5_N189_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_7_N189_PULSESHAPING (.ZN (N189), .A1 (XNOR_1_6_N189_PULSESHAPING_OUT), .A2 (GND));

      wire XNOR_1_1_N195_PULSESHAPING_OUT, XNOR_1_2_N195_PULSESHAPING_OUT, XNOR_1_3_N195_PULSESHAPING_OUT, XNOR_1_4_N195_PULSESHAPING_OUT, XNOR_1_5_N195_PULSESHAPING_OUT, XNOR_1_6_N195_PULSESHAPING_OUT;
      NOR2_X1 XNOR_1_1_N195_PULSESHAPING (.ZN (XNOR_1_1_N195_PULSESHAPING_OUT), .A1 (N195_PWL), .A2 (GND));
      NOR2_X1 XNOR_1_2_N195_PULSESHAPING (.ZN (XNOR_1_2_N195_PULSESHAPING_OUT), .A1 (XNOR_1_1_N195_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_3_N195_PULSESHAPING (.ZN (XNOR_1_3_N195_PULSESHAPING_OUT), .A1 (XNOR_1_2_N195_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_4_N195_PULSESHAPING (.ZN (XNOR_1_4_N195_PULSESHAPING_OUT), .A1 (XNOR_1_3_N195_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_5_N195_PULSESHAPING (.ZN (XNOR_1_5_N195_PULSESHAPING_OUT), .A1 (XNOR_1_4_N195_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_6_N195_PULSESHAPING (.ZN (XNOR_1_6_N195_PULSESHAPING_OUT), .A1 (XNOR_1_5_N195_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_7_N195_PULSESHAPING (.ZN (N195), .A1 (XNOR_1_6_N195_PULSESHAPING_OUT), .A2 (GND));

      wire XNOR_1_1_N201_PULSESHAPING_OUT, XNOR_1_2_N201_PULSESHAPING_OUT, XNOR_1_3_N201_PULSESHAPING_OUT, XNOR_1_4_N201_PULSESHAPING_OUT, XNOR_1_5_N201_PULSESHAPING_OUT, XNOR_1_6_N201_PULSESHAPING_OUT;
      NOR2_X1 XNOR_1_1_N201_PULSESHAPING (.ZN (XNOR_1_1_N201_PULSESHAPING_OUT), .A1 (N201_PWL), .A2 (GND));
      NOR2_X1 XNOR_1_2_N201_PULSESHAPING (.ZN (XNOR_1_2_N201_PULSESHAPING_OUT), .A1 (XNOR_1_1_N201_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_3_N201_PULSESHAPING (.ZN (XNOR_1_3_N201_PULSESHAPING_OUT), .A1 (XNOR_1_2_N201_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_4_N201_PULSESHAPING (.ZN (XNOR_1_4_N201_PULSESHAPING_OUT), .A1 (XNOR_1_3_N201_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_5_N201_PULSESHAPING (.ZN (XNOR_1_5_N201_PULSESHAPING_OUT), .A1 (XNOR_1_4_N201_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_6_N201_PULSESHAPING (.ZN (XNOR_1_6_N201_PULSESHAPING_OUT), .A1 (XNOR_1_5_N201_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_7_N201_PULSESHAPING (.ZN (N201), .A1 (XNOR_1_6_N201_PULSESHAPING_OUT), .A2 (GND));

      wire XNOR_1_1_N207_PULSESHAPING_OUT, XNOR_1_2_N207_PULSESHAPING_OUT, XNOR_1_3_N207_PULSESHAPING_OUT, XNOR_1_4_N207_PULSESHAPING_OUT, XNOR_1_5_N207_PULSESHAPING_OUT, XNOR_1_6_N207_PULSESHAPING_OUT;
      NOR2_X1 XNOR_1_1_N207_PULSESHAPING (.ZN (XNOR_1_1_N207_PULSESHAPING_OUT), .A1 (N207_PWL), .A2 (GND));
      NOR2_X1 XNOR_1_2_N207_PULSESHAPING (.ZN (XNOR_1_2_N207_PULSESHAPING_OUT), .A1 (XNOR_1_1_N207_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_3_N207_PULSESHAPING (.ZN (XNOR_1_3_N207_PULSESHAPING_OUT), .A1 (XNOR_1_2_N207_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_4_N207_PULSESHAPING (.ZN (XNOR_1_4_N207_PULSESHAPING_OUT), .A1 (XNOR_1_3_N207_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_5_N207_PULSESHAPING (.ZN (XNOR_1_5_N207_PULSESHAPING_OUT), .A1 (XNOR_1_4_N207_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_6_N207_PULSESHAPING (.ZN (XNOR_1_6_N207_PULSESHAPING_OUT), .A1 (XNOR_1_5_N207_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_7_N207_PULSESHAPING (.ZN (N207), .A1 (XNOR_1_6_N207_PULSESHAPING_OUT), .A2 (GND));

      wire XNOR_1_1_N210_PULSESHAPING_OUT, XNOR_1_2_N210_PULSESHAPING_OUT, XNOR_1_3_N210_PULSESHAPING_OUT, XNOR_1_4_N210_PULSESHAPING_OUT, XNOR_1_5_N210_PULSESHAPING_OUT, XNOR_1_6_N210_PULSESHAPING_OUT;
      NOR2_X1 XNOR_1_1_N210_PULSESHAPING (.ZN (XNOR_1_1_N210_PULSESHAPING_OUT), .A1 (N210_PWL), .A2 (GND));
      NOR2_X1 XNOR_1_2_N210_PULSESHAPING (.ZN (XNOR_1_2_N210_PULSESHAPING_OUT), .A1 (XNOR_1_1_N210_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_3_N210_PULSESHAPING (.ZN (XNOR_1_3_N210_PULSESHAPING_OUT), .A1 (XNOR_1_2_N210_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_4_N210_PULSESHAPING (.ZN (XNOR_1_4_N210_PULSESHAPING_OUT), .A1 (XNOR_1_3_N210_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_5_N210_PULSESHAPING (.ZN (XNOR_1_5_N210_PULSESHAPING_OUT), .A1 (XNOR_1_4_N210_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_6_N210_PULSESHAPING (.ZN (XNOR_1_6_N210_PULSESHAPING_OUT), .A1 (XNOR_1_5_N210_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_7_N210_PULSESHAPING (.ZN (N210), .A1 (XNOR_1_6_N210_PULSESHAPING_OUT), .A2 (GND));

      wire XNOR_1_1_N219_PULSESHAPING_OUT, XNOR_1_2_N219_PULSESHAPING_OUT, XNOR_1_3_N219_PULSESHAPING_OUT, XNOR_1_4_N219_PULSESHAPING_OUT, XNOR_1_5_N219_PULSESHAPING_OUT, XNOR_1_6_N219_PULSESHAPING_OUT;
      NOR2_X1 XNOR_1_1_N219_PULSESHAPING (.ZN (XNOR_1_1_N219_PULSESHAPING_OUT), .A1 (N219_PWL), .A2 (GND));
      NOR2_X1 XNOR_1_2_N219_PULSESHAPING (.ZN (XNOR_1_2_N219_PULSESHAPING_OUT), .A1 (XNOR_1_1_N219_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_3_N219_PULSESHAPING (.ZN (XNOR_1_3_N219_PULSESHAPING_OUT), .A1 (XNOR_1_2_N219_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_4_N219_PULSESHAPING (.ZN (XNOR_1_4_N219_PULSESHAPING_OUT), .A1 (XNOR_1_3_N219_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_5_N219_PULSESHAPING (.ZN (XNOR_1_5_N219_PULSESHAPING_OUT), .A1 (XNOR_1_4_N219_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_6_N219_PULSESHAPING (.ZN (XNOR_1_6_N219_PULSESHAPING_OUT), .A1 (XNOR_1_5_N219_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_7_N219_PULSESHAPING (.ZN (N219), .A1 (XNOR_1_6_N219_PULSESHAPING_OUT), .A2 (GND));

      wire XNOR_1_1_N228_PULSESHAPING_OUT, XNOR_1_2_N228_PULSESHAPING_OUT, XNOR_1_3_N228_PULSESHAPING_OUT, XNOR_1_4_N228_PULSESHAPING_OUT, XNOR_1_5_N228_PULSESHAPING_OUT, XNOR_1_6_N228_PULSESHAPING_OUT;
      NOR2_X1 XNOR_1_1_N228_PULSESHAPING (.ZN (XNOR_1_1_N228_PULSESHAPING_OUT), .A1 (N228_PWL), .A2 (GND));
      NOR2_X1 XNOR_1_2_N228_PULSESHAPING (.ZN (XNOR_1_2_N228_PULSESHAPING_OUT), .A1 (XNOR_1_1_N228_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_3_N228_PULSESHAPING (.ZN (XNOR_1_3_N228_PULSESHAPING_OUT), .A1 (XNOR_1_2_N228_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_4_N228_PULSESHAPING (.ZN (XNOR_1_4_N228_PULSESHAPING_OUT), .A1 (XNOR_1_3_N228_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_5_N228_PULSESHAPING (.ZN (XNOR_1_5_N228_PULSESHAPING_OUT), .A1 (XNOR_1_4_N228_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_6_N228_PULSESHAPING (.ZN (XNOR_1_6_N228_PULSESHAPING_OUT), .A1 (XNOR_1_5_N228_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_7_N228_PULSESHAPING (.ZN (N228), .A1 (XNOR_1_6_N228_PULSESHAPING_OUT), .A2 (GND));

      wire XNOR_1_1_N237_PULSESHAPING_OUT, XNOR_1_2_N237_PULSESHAPING_OUT, XNOR_1_3_N237_PULSESHAPING_OUT, XNOR_1_4_N237_PULSESHAPING_OUT, XNOR_1_5_N237_PULSESHAPING_OUT, XNOR_1_6_N237_PULSESHAPING_OUT;
      NOR2_X1 XNOR_1_1_N237_PULSESHAPING (.ZN (XNOR_1_1_N237_PULSESHAPING_OUT), .A1 (N237_PWL), .A2 (GND));
      NOR2_X1 XNOR_1_2_N237_PULSESHAPING (.ZN (XNOR_1_2_N237_PULSESHAPING_OUT), .A1 (XNOR_1_1_N237_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_3_N237_PULSESHAPING (.ZN (XNOR_1_3_N237_PULSESHAPING_OUT), .A1 (XNOR_1_2_N237_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_4_N237_PULSESHAPING (.ZN (XNOR_1_4_N237_PULSESHAPING_OUT), .A1 (XNOR_1_3_N237_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_5_N237_PULSESHAPING (.ZN (XNOR_1_5_N237_PULSESHAPING_OUT), .A1 (XNOR_1_4_N237_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_6_N237_PULSESHAPING (.ZN (XNOR_1_6_N237_PULSESHAPING_OUT), .A1 (XNOR_1_5_N237_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_7_N237_PULSESHAPING (.ZN (N237), .A1 (XNOR_1_6_N237_PULSESHAPING_OUT), .A2 (GND));

      wire XNOR_1_1_N246_PULSESHAPING_OUT, XNOR_1_2_N246_PULSESHAPING_OUT, XNOR_1_3_N246_PULSESHAPING_OUT, XNOR_1_4_N246_PULSESHAPING_OUT, XNOR_1_5_N246_PULSESHAPING_OUT, XNOR_1_6_N246_PULSESHAPING_OUT;
      NOR2_X1 XNOR_1_1_N246_PULSESHAPING (.ZN (XNOR_1_1_N246_PULSESHAPING_OUT), .A1 (N246_PWL), .A2 (GND));
      NOR2_X1 XNOR_1_2_N246_PULSESHAPING (.ZN (XNOR_1_2_N246_PULSESHAPING_OUT), .A1 (XNOR_1_1_N246_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_3_N246_PULSESHAPING (.ZN (XNOR_1_3_N246_PULSESHAPING_OUT), .A1 (XNOR_1_2_N246_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_4_N246_PULSESHAPING (.ZN (XNOR_1_4_N246_PULSESHAPING_OUT), .A1 (XNOR_1_3_N246_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_5_N246_PULSESHAPING (.ZN (XNOR_1_5_N246_PULSESHAPING_OUT), .A1 (XNOR_1_4_N246_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_6_N246_PULSESHAPING (.ZN (XNOR_1_6_N246_PULSESHAPING_OUT), .A1 (XNOR_1_5_N246_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_7_N246_PULSESHAPING (.ZN (N246), .A1 (XNOR_1_6_N246_PULSESHAPING_OUT), .A2 (GND));

      wire XNOR_1_1_N255_PULSESHAPING_OUT, XNOR_1_2_N255_PULSESHAPING_OUT, XNOR_1_3_N255_PULSESHAPING_OUT, XNOR_1_4_N255_PULSESHAPING_OUT, XNOR_1_5_N255_PULSESHAPING_OUT, XNOR_1_6_N255_PULSESHAPING_OUT;
      NOR2_X1 XNOR_1_1_N255_PULSESHAPING (.ZN (XNOR_1_1_N255_PULSESHAPING_OUT), .A1 (N255_PWL), .A2 (GND));
      NOR2_X1 XNOR_1_2_N255_PULSESHAPING (.ZN (XNOR_1_2_N255_PULSESHAPING_OUT), .A1 (XNOR_1_1_N255_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_3_N255_PULSESHAPING (.ZN (XNOR_1_3_N255_PULSESHAPING_OUT), .A1 (XNOR_1_2_N255_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_4_N255_PULSESHAPING (.ZN (XNOR_1_4_N255_PULSESHAPING_OUT), .A1 (XNOR_1_3_N255_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_5_N255_PULSESHAPING (.ZN (XNOR_1_5_N255_PULSESHAPING_OUT), .A1 (XNOR_1_4_N255_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_6_N255_PULSESHAPING (.ZN (XNOR_1_6_N255_PULSESHAPING_OUT), .A1 (XNOR_1_5_N255_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_7_N255_PULSESHAPING (.ZN (N255), .A1 (XNOR_1_6_N255_PULSESHAPING_OUT), .A2 (GND));

      wire XNOR_1_1_N259_PULSESHAPING_OUT, XNOR_1_2_N259_PULSESHAPING_OUT, XNOR_1_3_N259_PULSESHAPING_OUT, XNOR_1_4_N259_PULSESHAPING_OUT, XNOR_1_5_N259_PULSESHAPING_OUT, XNOR_1_6_N259_PULSESHAPING_OUT;
      NOR2_X1 XNOR_1_1_N259_PULSESHAPING (.ZN (XNOR_1_1_N259_PULSESHAPING_OUT), .A1 (N259_PWL), .A2 (GND));
      NOR2_X1 XNOR_1_2_N259_PULSESHAPING (.ZN (XNOR_1_2_N259_PULSESHAPING_OUT), .A1 (XNOR_1_1_N259_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_3_N259_PULSESHAPING (.ZN (XNOR_1_3_N259_PULSESHAPING_OUT), .A1 (XNOR_1_2_N259_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_4_N259_PULSESHAPING (.ZN (XNOR_1_4_N259_PULSESHAPING_OUT), .A1 (XNOR_1_3_N259_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_5_N259_PULSESHAPING (.ZN (XNOR_1_5_N259_PULSESHAPING_OUT), .A1 (XNOR_1_4_N259_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_6_N259_PULSESHAPING (.ZN (XNOR_1_6_N259_PULSESHAPING_OUT), .A1 (XNOR_1_5_N259_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_7_N259_PULSESHAPING (.ZN (N259), .A1 (XNOR_1_6_N259_PULSESHAPING_OUT), .A2 (GND));

      wire XNOR_1_1_N260_PULSESHAPING_OUT, XNOR_1_2_N260_PULSESHAPING_OUT, XNOR_1_3_N260_PULSESHAPING_OUT, XNOR_1_4_N260_PULSESHAPING_OUT, XNOR_1_5_N260_PULSESHAPING_OUT, XNOR_1_6_N260_PULSESHAPING_OUT;
      NOR2_X1 XNOR_1_1_N260_PULSESHAPING (.ZN (XNOR_1_1_N260_PULSESHAPING_OUT), .A1 (N260_PWL), .A2 (GND));
      NOR2_X1 XNOR_1_2_N260_PULSESHAPING (.ZN (XNOR_1_2_N260_PULSESHAPING_OUT), .A1 (XNOR_1_1_N260_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_3_N260_PULSESHAPING (.ZN (XNOR_1_3_N260_PULSESHAPING_OUT), .A1 (XNOR_1_2_N260_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_4_N260_PULSESHAPING (.ZN (XNOR_1_4_N260_PULSESHAPING_OUT), .A1 (XNOR_1_3_N260_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_5_N260_PULSESHAPING (.ZN (XNOR_1_5_N260_PULSESHAPING_OUT), .A1 (XNOR_1_4_N260_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_6_N260_PULSESHAPING (.ZN (XNOR_1_6_N260_PULSESHAPING_OUT), .A1 (XNOR_1_5_N260_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_7_N260_PULSESHAPING (.ZN (N260), .A1 (XNOR_1_6_N260_PULSESHAPING_OUT), .A2 (GND));

      wire XNOR_1_1_N261_PULSESHAPING_OUT, XNOR_1_2_N261_PULSESHAPING_OUT, XNOR_1_3_N261_PULSESHAPING_OUT, XNOR_1_4_N261_PULSESHAPING_OUT, XNOR_1_5_N261_PULSESHAPING_OUT, XNOR_1_6_N261_PULSESHAPING_OUT;
      NOR2_X1 XNOR_1_1_N261_PULSESHAPING (.ZN (XNOR_1_1_N261_PULSESHAPING_OUT), .A1 (N261_PWL), .A2 (GND));
      NOR2_X1 XNOR_1_2_N261_PULSESHAPING (.ZN (XNOR_1_2_N261_PULSESHAPING_OUT), .A1 (XNOR_1_1_N261_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_3_N261_PULSESHAPING (.ZN (XNOR_1_3_N261_PULSESHAPING_OUT), .A1 (XNOR_1_2_N261_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_4_N261_PULSESHAPING (.ZN (XNOR_1_4_N261_PULSESHAPING_OUT), .A1 (XNOR_1_3_N261_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_5_N261_PULSESHAPING (.ZN (XNOR_1_5_N261_PULSESHAPING_OUT), .A1 (XNOR_1_4_N261_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_6_N261_PULSESHAPING (.ZN (XNOR_1_6_N261_PULSESHAPING_OUT), .A1 (XNOR_1_5_N261_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_7_N261_PULSESHAPING (.ZN (N261), .A1 (XNOR_1_6_N261_PULSESHAPING_OUT), .A2 (GND));

      wire XNOR_1_1_N267_PULSESHAPING_OUT, XNOR_1_2_N267_PULSESHAPING_OUT, XNOR_1_3_N267_PULSESHAPING_OUT, XNOR_1_4_N267_PULSESHAPING_OUT, XNOR_1_5_N267_PULSESHAPING_OUT, XNOR_1_6_N267_PULSESHAPING_OUT;
      NOR2_X1 XNOR_1_1_N267_PULSESHAPING (.ZN (XNOR_1_1_N267_PULSESHAPING_OUT), .A1 (N267_PWL), .A2 (GND));
      NOR2_X1 XNOR_1_2_N267_PULSESHAPING (.ZN (XNOR_1_2_N267_PULSESHAPING_OUT), .A1 (XNOR_1_1_N267_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_3_N267_PULSESHAPING (.ZN (XNOR_1_3_N267_PULSESHAPING_OUT), .A1 (XNOR_1_2_N267_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_4_N267_PULSESHAPING (.ZN (XNOR_1_4_N267_PULSESHAPING_OUT), .A1 (XNOR_1_3_N267_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_5_N267_PULSESHAPING (.ZN (XNOR_1_5_N267_PULSESHAPING_OUT), .A1 (XNOR_1_4_N267_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_6_N267_PULSESHAPING (.ZN (XNOR_1_6_N267_PULSESHAPING_OUT), .A1 (XNOR_1_5_N267_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_7_N267_PULSESHAPING (.ZN (N267), .A1 (XNOR_1_6_N267_PULSESHAPING_OUT), .A2 (GND));

      wire XNOR_1_1_N268_PULSESHAPING_OUT, XNOR_1_2_N268_PULSESHAPING_OUT, XNOR_1_3_N268_PULSESHAPING_OUT, XNOR_1_4_N268_PULSESHAPING_OUT, XNOR_1_5_N268_PULSESHAPING_OUT, XNOR_1_6_N268_PULSESHAPING_OUT;
      NOR2_X1 XNOR_1_1_N268_PULSESHAPING (.ZN (XNOR_1_1_N268_PULSESHAPING_OUT), .A1 (N268_PWL), .A2 (GND));
      NOR2_X1 XNOR_1_2_N268_PULSESHAPING (.ZN (XNOR_1_2_N268_PULSESHAPING_OUT), .A1 (XNOR_1_1_N268_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_3_N268_PULSESHAPING (.ZN (XNOR_1_3_N268_PULSESHAPING_OUT), .A1 (XNOR_1_2_N268_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_4_N268_PULSESHAPING (.ZN (XNOR_1_4_N268_PULSESHAPING_OUT), .A1 (XNOR_1_3_N268_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_5_N268_PULSESHAPING (.ZN (XNOR_1_5_N268_PULSESHAPING_OUT), .A1 (XNOR_1_4_N268_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_6_N268_PULSESHAPING (.ZN (XNOR_1_6_N268_PULSESHAPING_OUT), .A1 (XNOR_1_5_N268_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_7_N268_PULSESHAPING (.ZN (N268), .A1 (XNOR_1_6_N268_PULSESHAPING_OUT), .A2 (GND));



      wire XNOR_1_1_NUM1_OUT, XNOR_1_2_NUM1_OUT, XNOR_1_3_NUM1_OUT;
      NOR2_X1 XNOR_1_1_NUM1 (.ZN (XNOR_1_1_NUM1_OUT), .A1 (N1), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM1 (.ZN (XNOR_1_2_NUM1_OUT), .A1 (GND), .A2 (N8));
      NOR2_X1 XNOR_1_3_NUM1 (.ZN (XNOR_1_3_NUM1_OUT), .A1 (XNOR_1_1_NUM1_OUT), .A2 (XNOR_1_2_NUM1_OUT));

      wire XNOR_2_1_NUM1_OUT, XNOR_2_2_NUM1_OUT, XNOR_2_3_NUM1_OUT;
      NOR2_X1 XNOR_2_1_NUM1 (.ZN (XNOR_2_1_NUM1_OUT), .A1 (N13), .A2 (GND));
      NOR2_X1 XNOR_2_2_NUM1 (.ZN (XNOR_2_2_NUM1_OUT), .A1 (GND), .A2 (N17));
      NOR2_X1 XNOR_2_3_NUM1 (.ZN (XNOR_2_3_NUM1_OUT), .A1 (XNOR_2_1_NUM1_OUT), .A2 (XNOR_2_2_NUM1_OUT));

      wire XNOR_3_1_NUM1_OUT, XNOR_3_2_NUM1_OUT, XNOR_3_3_NUM1_OUT;
      NOR2_X1 XNOR_3_1_NUM1 (.ZN (XNOR_3_1_NUM1_OUT), .A1 (XNOR_1_3_NUM1_OUT), .A2 (GND));
      NOR2_X1 XNOR_3_2_NUM1 (.ZN (XNOR_3_2_NUM1_OUT), .A1 (GND), .A2 (XNOR_2_3_NUM1_OUT));
      NOR2_X1 XNOR_3_3_NUM1 (.ZN (XNOR_3_3_NUM1_OUT), .A1 (XNOR_3_1_NUM1_OUT), .A2 (XNOR_3_2_NUM1_OUT));

      NOR2_X1 XNOR_4_1_NUM1 (.ZN (N269), .A1 (XNOR_3_3_NUM1_OUT), .A2 (GND));
      wire XNOR_1_1_NUM2_OUT, XNOR_1_2_NUM2_OUT, XNOR_1_3_NUM2_OUT;
      NOR2_X1 XNOR_1_1_NUM2 (.ZN (XNOR_1_1_NUM2_OUT), .A1 (N1), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM2 (.ZN (XNOR_1_2_NUM2_OUT), .A1 (GND), .A2 (N26));
      NOR2_X1 XNOR_1_3_NUM2 (.ZN (XNOR_1_3_NUM2_OUT), .A1 (XNOR_1_1_NUM2_OUT), .A2 (XNOR_1_2_NUM2_OUT));

      wire XNOR_2_1_NUM2_OUT, XNOR_2_2_NUM2_OUT, XNOR_2_3_NUM2_OUT;
      NOR2_X1 XNOR_2_1_NUM2 (.ZN (XNOR_2_1_NUM2_OUT), .A1 (N13), .A2 (GND));
      NOR2_X1 XNOR_2_2_NUM2 (.ZN (XNOR_2_2_NUM2_OUT), .A1 (GND), .A2 (N17));
      NOR2_X1 XNOR_2_3_NUM2 (.ZN (XNOR_2_3_NUM2_OUT), .A1 (XNOR_2_1_NUM2_OUT), .A2 (XNOR_2_2_NUM2_OUT));

      wire XNOR_3_1_NUM2_OUT, XNOR_3_2_NUM2_OUT, XNOR_3_3_NUM2_OUT;
      NOR2_X1 XNOR_3_1_NUM2 (.ZN (XNOR_3_1_NUM2_OUT), .A1 (XNOR_1_3_NUM2_OUT), .A2 (GND));
      NOR2_X1 XNOR_3_2_NUM2 (.ZN (XNOR_3_2_NUM2_OUT), .A1 (GND), .A2 (XNOR_2_3_NUM2_OUT));
      NOR2_X1 XNOR_3_3_NUM2 (.ZN (XNOR_3_3_NUM2_OUT), .A1 (XNOR_3_1_NUM2_OUT), .A2 (XNOR_3_2_NUM2_OUT));

      NOR2_X1 XNOR_4_1_NUM2 (.ZN (N270), .A1 (XNOR_3_3_NUM2_OUT), .A2 (GND));
      wire XNOR_1_1_NUM3_OUT, XNOR_1_2_NUM3_OUT, XNOR_1_3_NUM3_OUT;
      NOR2_X1 XNOR_1_1_NUM3 (.ZN (XNOR_1_1_NUM3_OUT), .A1 (N29), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM3 (.ZN (XNOR_1_2_NUM3_OUT), .A1 (GND), .A2 (N36));
      NOR2_X1 XNOR_1_3_NUM3 (.ZN (XNOR_1_3_NUM3_OUT), .A1 (XNOR_1_1_NUM3_OUT), .A2 (XNOR_1_2_NUM3_OUT));

      wire XNOR_2_1_NUM3_OUT, XNOR_2_2_NUM3_OUT;
      NOR2_X1 XNOR_2_1_NUM3 (.ZN (XNOR_2_1_NUM3_OUT), .A1 (N42), .A2 (GND));
      NOR2_X1 XNOR_2_2_NUM3 (.ZN (XNOR_2_2_NUM3_OUT), .A1 (GND), .A2 (XNOR_1_3_NUM3_OUT));
      NOR2_X1 XNOR_2_3_NUM3 (.ZN (N273), .A1 (XNOR_2_1_NUM3_OUT), .A2 (XNOR_2_2_NUM3_OUT));
      wire XNOR_1_1_NUM4_OUT, XNOR_1_2_NUM4_OUT, XNOR_1_3_NUM4_OUT;
      NOR2_X1 XNOR_1_1_NUM4 (.ZN (XNOR_1_1_NUM4_OUT), .A1 (N1), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM4 (.ZN (XNOR_1_2_NUM4_OUT), .A1 (GND), .A2 (N26));
      NOR2_X1 XNOR_1_3_NUM4 (.ZN (XNOR_1_3_NUM4_OUT), .A1 (XNOR_1_1_NUM4_OUT), .A2 (XNOR_1_2_NUM4_OUT));

      wire XNOR_2_1_NUM4_OUT, XNOR_2_2_NUM4_OUT;
      NOR2_X1 XNOR_2_1_NUM4 (.ZN (XNOR_2_1_NUM4_OUT), .A1 (N51), .A2 (GND));
      NOR2_X1 XNOR_2_2_NUM4 (.ZN (XNOR_2_2_NUM4_OUT), .A1 (GND), .A2 (XNOR_1_3_NUM4_OUT));
      NOR2_X1 XNOR_2_3_NUM4 (.ZN (N276), .A1 (XNOR_2_1_NUM4_OUT), .A2 (XNOR_2_2_NUM4_OUT));
      wire XNOR_1_1_NUM5_OUT, XNOR_1_2_NUM5_OUT, XNOR_1_3_NUM5_OUT;
      NOR2_X1 XNOR_1_1_NUM5 (.ZN (XNOR_1_1_NUM5_OUT), .A1 (N1), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM5 (.ZN (XNOR_1_2_NUM5_OUT), .A1 (GND), .A2 (N8));
      NOR2_X1 XNOR_1_3_NUM5 (.ZN (XNOR_1_3_NUM5_OUT), .A1 (XNOR_1_1_NUM5_OUT), .A2 (XNOR_1_2_NUM5_OUT));

      wire XNOR_2_1_NUM5_OUT, XNOR_2_2_NUM5_OUT, XNOR_2_3_NUM5_OUT;
      NOR2_X1 XNOR_2_1_NUM5 (.ZN (XNOR_2_1_NUM5_OUT), .A1 (N51), .A2 (GND));
      NOR2_X1 XNOR_2_2_NUM5 (.ZN (XNOR_2_2_NUM5_OUT), .A1 (GND), .A2 (N17));
      NOR2_X1 XNOR_2_3_NUM5 (.ZN (XNOR_2_3_NUM5_OUT), .A1 (XNOR_2_1_NUM5_OUT), .A2 (XNOR_2_2_NUM5_OUT));

      wire XNOR_3_1_NUM5_OUT, XNOR_3_2_NUM5_OUT, XNOR_3_3_NUM5_OUT;
      NOR2_X1 XNOR_3_1_NUM5 (.ZN (XNOR_3_1_NUM5_OUT), .A1 (XNOR_1_3_NUM5_OUT), .A2 (GND));
      NOR2_X1 XNOR_3_2_NUM5 (.ZN (XNOR_3_2_NUM5_OUT), .A1 (GND), .A2 (XNOR_2_3_NUM5_OUT));
      NOR2_X1 XNOR_3_3_NUM5 (.ZN (XNOR_3_3_NUM5_OUT), .A1 (XNOR_3_1_NUM5_OUT), .A2 (XNOR_3_2_NUM5_OUT));

      NOR2_X1 XNOR_4_1_NUM5 (.ZN (N279), .A1 (XNOR_3_3_NUM5_OUT), .A2 (GND));
      wire XNOR_1_1_NUM6_OUT, XNOR_1_2_NUM6_OUT, XNOR_1_3_NUM6_OUT;
      NOR2_X1 XNOR_1_1_NUM6 (.ZN (XNOR_1_1_NUM6_OUT), .A1 (N1), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM6 (.ZN (XNOR_1_2_NUM6_OUT), .A1 (GND), .A2 (N8));
      NOR2_X1 XNOR_1_3_NUM6 (.ZN (XNOR_1_3_NUM6_OUT), .A1 (XNOR_1_1_NUM6_OUT), .A2 (XNOR_1_2_NUM6_OUT));

      wire XNOR_2_1_NUM6_OUT, XNOR_2_2_NUM6_OUT, XNOR_2_3_NUM6_OUT;
      NOR2_X1 XNOR_2_1_NUM6 (.ZN (XNOR_2_1_NUM6_OUT), .A1 (N13), .A2 (GND));
      NOR2_X1 XNOR_2_2_NUM6 (.ZN (XNOR_2_2_NUM6_OUT), .A1 (GND), .A2 (N55));
      NOR2_X1 XNOR_2_3_NUM6 (.ZN (XNOR_2_3_NUM6_OUT), .A1 (XNOR_2_1_NUM6_OUT), .A2 (XNOR_2_2_NUM6_OUT));

      wire XNOR_3_1_NUM6_OUT, XNOR_3_2_NUM6_OUT, XNOR_3_3_NUM6_OUT;
      NOR2_X1 XNOR_3_1_NUM6 (.ZN (XNOR_3_1_NUM6_OUT), .A1 (XNOR_1_3_NUM6_OUT), .A2 (GND));
      NOR2_X1 XNOR_3_2_NUM6 (.ZN (XNOR_3_2_NUM6_OUT), .A1 (GND), .A2 (XNOR_2_3_NUM6_OUT));
      NOR2_X1 XNOR_3_3_NUM6 (.ZN (XNOR_3_3_NUM6_OUT), .A1 (XNOR_3_1_NUM6_OUT), .A2 (XNOR_3_2_NUM6_OUT));

      NOR2_X1 XNOR_4_1_NUM6 (.ZN (N280), .A1 (XNOR_3_3_NUM6_OUT), .A2 (GND));
      wire XNOR_1_1_NUM7_OUT, XNOR_1_2_NUM7_OUT, XNOR_1_3_NUM7_OUT;
      NOR2_X1 XNOR_1_1_NUM7 (.ZN (XNOR_1_1_NUM7_OUT), .A1 (N59), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM7 (.ZN (XNOR_1_2_NUM7_OUT), .A1 (GND), .A2 (N42));
      NOR2_X1 XNOR_1_3_NUM7 (.ZN (XNOR_1_3_NUM7_OUT), .A1 (XNOR_1_1_NUM7_OUT), .A2 (XNOR_1_2_NUM7_OUT));

      wire XNOR_2_1_NUM7_OUT, XNOR_2_2_NUM7_OUT, XNOR_2_3_NUM7_OUT;
      NOR2_X1 XNOR_2_1_NUM7 (.ZN (XNOR_2_1_NUM7_OUT), .A1 (N68), .A2 (GND));
      NOR2_X1 XNOR_2_2_NUM7 (.ZN (XNOR_2_2_NUM7_OUT), .A1 (GND), .A2 (N72));
      NOR2_X1 XNOR_2_3_NUM7 (.ZN (XNOR_2_3_NUM7_OUT), .A1 (XNOR_2_1_NUM7_OUT), .A2 (XNOR_2_2_NUM7_OUT));

      wire XNOR_3_1_NUM7_OUT, XNOR_3_2_NUM7_OUT, XNOR_3_3_NUM7_OUT;
      NOR2_X1 XNOR_3_1_NUM7 (.ZN (XNOR_3_1_NUM7_OUT), .A1 (XNOR_1_3_NUM7_OUT), .A2 (GND));
      NOR2_X1 XNOR_3_2_NUM7 (.ZN (XNOR_3_2_NUM7_OUT), .A1 (GND), .A2 (XNOR_2_3_NUM7_OUT));
      NOR2_X1 XNOR_3_3_NUM7 (.ZN (XNOR_3_3_NUM7_OUT), .A1 (XNOR_3_1_NUM7_OUT), .A2 (XNOR_3_2_NUM7_OUT));

      NOR2_X1 XNOR_4_1_NUM7 (.ZN (N284), .A1 (XNOR_3_3_NUM7_OUT), .A2 (GND));
      wire XNOR_1_1_NUM8_OUT, XNOR_1_2_NUM8_OUT, XNOR_1_3_NUM8_OUT;
      NOR2_X1 XNOR_1_1_NUM8 (.ZN (XNOR_1_1_NUM8_OUT), .A1 (N29), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM8 (.ZN (XNOR_1_2_NUM8_OUT), .A1 (GND), .A2 (N68));
      NOR2_X1 XNOR_1_3_NUM8 (.ZN (XNOR_1_3_NUM8_OUT), .A1 (XNOR_1_1_NUM8_OUT), .A2 (XNOR_1_2_NUM8_OUT));
      NOR2_X1 XNOR_1_4_NUM8 (.ZN (N285), .A1 (XNOR_1_3_NUM8_OUT), .A2 (GND));
      wire XNOR_1_1_NUM9_OUT, XNOR_1_2_NUM9_OUT, XNOR_1_3_NUM9_OUT;
      NOR2_X1 XNOR_1_1_NUM9 (.ZN (XNOR_1_1_NUM9_OUT), .A1 (N59), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM9 (.ZN (XNOR_1_2_NUM9_OUT), .A1 (GND), .A2 (N68));
      NOR2_X1 XNOR_1_3_NUM9 (.ZN (XNOR_1_3_NUM9_OUT), .A1 (XNOR_1_1_NUM9_OUT), .A2 (XNOR_1_2_NUM9_OUT));

      wire XNOR_2_1_NUM9_OUT, XNOR_2_2_NUM9_OUT, XNOR_2_3_NUM9_OUT;
      NOR2_X1 XNOR_2_1_NUM9 (.ZN (XNOR_2_1_NUM9_OUT), .A1 (N74), .A2 (GND));
      NOR2_X1 XNOR_2_2_NUM9 (.ZN (XNOR_2_2_NUM9_OUT), .A1 (GND), .A2 (XNOR_1_3_NUM9_OUT));
      NOR2_X1 XNOR_2_3_NUM9 (.ZN (XNOR_2_3_NUM9_OUT), .A1 (XNOR_2_1_NUM9_OUT), .A2 (XNOR_2_2_NUM9_OUT));

      NOR2_X1 XNOR_3_1_NUM9 (.ZN (N286), .A1 (XNOR_2_3_NUM9_OUT), .A2 (GND));
      wire XNOR_1_1_NUM10_OUT, XNOR_1_2_NUM10_OUT, XNOR_1_3_NUM10_OUT;
      NOR2_X1 XNOR_1_1_NUM10 (.ZN (XNOR_1_1_NUM10_OUT), .A1 (N29), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM10 (.ZN (XNOR_1_2_NUM10_OUT), .A1 (GND), .A2 (N75));
      NOR2_X1 XNOR_1_3_NUM10 (.ZN (XNOR_1_3_NUM10_OUT), .A1 (XNOR_1_1_NUM10_OUT), .A2 (XNOR_1_2_NUM10_OUT));

      wire XNOR_2_1_NUM10_OUT, XNOR_2_2_NUM10_OUT;
      NOR2_X1 XNOR_2_1_NUM10 (.ZN (XNOR_2_1_NUM10_OUT), .A1 (N80), .A2 (GND));
      NOR2_X1 XNOR_2_2_NUM10 (.ZN (XNOR_2_2_NUM10_OUT), .A1 (GND), .A2 (XNOR_1_3_NUM10_OUT));
      NOR2_X1 XNOR_2_3_NUM10 (.ZN (N287), .A1 (XNOR_2_1_NUM10_OUT), .A2 (XNOR_2_2_NUM10_OUT));
      wire XNOR_1_1_NUM11_OUT, XNOR_1_2_NUM11_OUT, XNOR_1_3_NUM11_OUT;
      NOR2_X1 XNOR_1_1_NUM11 (.ZN (XNOR_1_1_NUM11_OUT), .A1 (N29), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM11 (.ZN (XNOR_1_2_NUM11_OUT), .A1 (GND), .A2 (N75));
      NOR2_X1 XNOR_1_3_NUM11 (.ZN (XNOR_1_3_NUM11_OUT), .A1 (XNOR_1_1_NUM11_OUT), .A2 (XNOR_1_2_NUM11_OUT));

      wire XNOR_2_1_NUM11_OUT, XNOR_2_2_NUM11_OUT;
      NOR2_X1 XNOR_2_1_NUM11 (.ZN (XNOR_2_1_NUM11_OUT), .A1 (N42), .A2 (GND));
      NOR2_X1 XNOR_2_2_NUM11 (.ZN (XNOR_2_2_NUM11_OUT), .A1 (GND), .A2 (XNOR_1_3_NUM11_OUT));
      NOR2_X1 XNOR_2_3_NUM11 (.ZN (N290), .A1 (XNOR_2_1_NUM11_OUT), .A2 (XNOR_2_2_NUM11_OUT));
      wire XNOR_1_1_NUM12_OUT, XNOR_1_2_NUM12_OUT, XNOR_1_3_NUM12_OUT;
      NOR2_X1 XNOR_1_1_NUM12 (.ZN (XNOR_1_1_NUM12_OUT), .A1 (N29), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM12 (.ZN (XNOR_1_2_NUM12_OUT), .A1 (GND), .A2 (N36));
      NOR2_X1 XNOR_1_3_NUM12 (.ZN (XNOR_1_3_NUM12_OUT), .A1 (XNOR_1_1_NUM12_OUT), .A2 (XNOR_1_2_NUM12_OUT));

      wire XNOR_2_1_NUM12_OUT, XNOR_2_2_NUM12_OUT;
      NOR2_X1 XNOR_2_1_NUM12 (.ZN (XNOR_2_1_NUM12_OUT), .A1 (N80), .A2 (GND));
      NOR2_X1 XNOR_2_2_NUM12 (.ZN (XNOR_2_2_NUM12_OUT), .A1 (GND), .A2 (XNOR_1_3_NUM12_OUT));
      NOR2_X1 XNOR_2_3_NUM12 (.ZN (N291), .A1 (XNOR_2_1_NUM12_OUT), .A2 (XNOR_2_2_NUM12_OUT));
      wire XNOR_1_1_NUM13_OUT, XNOR_1_2_NUM13_OUT, XNOR_1_3_NUM13_OUT;
      NOR2_X1 XNOR_1_1_NUM13 (.ZN (XNOR_1_1_NUM13_OUT), .A1 (N29), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM13 (.ZN (XNOR_1_2_NUM13_OUT), .A1 (GND), .A2 (N36));
      NOR2_X1 XNOR_1_3_NUM13 (.ZN (XNOR_1_3_NUM13_OUT), .A1 (XNOR_1_1_NUM13_OUT), .A2 (XNOR_1_2_NUM13_OUT));

      wire XNOR_2_1_NUM13_OUT, XNOR_2_2_NUM13_OUT;
      NOR2_X1 XNOR_2_1_NUM13 (.ZN (XNOR_2_1_NUM13_OUT), .A1 (N42), .A2 (GND));
      NOR2_X1 XNOR_2_2_NUM13 (.ZN (XNOR_2_2_NUM13_OUT), .A1 (GND), .A2 (XNOR_1_3_NUM13_OUT));
      NOR2_X1 XNOR_2_3_NUM13 (.ZN (N292), .A1 (XNOR_2_1_NUM13_OUT), .A2 (XNOR_2_2_NUM13_OUT));
      wire XNOR_1_1_NUM14_OUT, XNOR_1_2_NUM14_OUT, XNOR_1_3_NUM14_OUT;
      NOR2_X1 XNOR_1_1_NUM14 (.ZN (XNOR_1_1_NUM14_OUT), .A1 (N59), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM14 (.ZN (XNOR_1_2_NUM14_OUT), .A1 (GND), .A2 (N75));
      NOR2_X1 XNOR_1_3_NUM14 (.ZN (XNOR_1_3_NUM14_OUT), .A1 (XNOR_1_1_NUM14_OUT), .A2 (XNOR_1_2_NUM14_OUT));

      wire XNOR_2_1_NUM14_OUT, XNOR_2_2_NUM14_OUT;
      NOR2_X1 XNOR_2_1_NUM14 (.ZN (XNOR_2_1_NUM14_OUT), .A1 (N80), .A2 (GND));
      NOR2_X1 XNOR_2_2_NUM14 (.ZN (XNOR_2_2_NUM14_OUT), .A1 (GND), .A2 (XNOR_1_3_NUM14_OUT));
      NOR2_X1 XNOR_2_3_NUM14 (.ZN (N293), .A1 (XNOR_2_1_NUM14_OUT), .A2 (XNOR_2_2_NUM14_OUT));
      wire XNOR_1_1_NUM15_OUT, XNOR_1_2_NUM15_OUT, XNOR_1_3_NUM15_OUT;
      NOR2_X1 XNOR_1_1_NUM15 (.ZN (XNOR_1_1_NUM15_OUT), .A1 (N59), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM15 (.ZN (XNOR_1_2_NUM15_OUT), .A1 (GND), .A2 (N75));
      NOR2_X1 XNOR_1_3_NUM15 (.ZN (XNOR_1_3_NUM15_OUT), .A1 (XNOR_1_1_NUM15_OUT), .A2 (XNOR_1_2_NUM15_OUT));

      wire XNOR_2_1_NUM15_OUT, XNOR_2_2_NUM15_OUT;
      NOR2_X1 XNOR_2_1_NUM15 (.ZN (XNOR_2_1_NUM15_OUT), .A1 (N42), .A2 (GND));
      NOR2_X1 XNOR_2_2_NUM15 (.ZN (XNOR_2_2_NUM15_OUT), .A1 (GND), .A2 (XNOR_1_3_NUM15_OUT));
      NOR2_X1 XNOR_2_3_NUM15 (.ZN (N294), .A1 (XNOR_2_1_NUM15_OUT), .A2 (XNOR_2_2_NUM15_OUT));
      wire XNOR_1_1_NUM16_OUT, XNOR_1_2_NUM16_OUT, XNOR_1_3_NUM16_OUT;
      NOR2_X1 XNOR_1_1_NUM16 (.ZN (XNOR_1_1_NUM16_OUT), .A1 (N59), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM16 (.ZN (XNOR_1_2_NUM16_OUT), .A1 (GND), .A2 (N36));
      NOR2_X1 XNOR_1_3_NUM16 (.ZN (XNOR_1_3_NUM16_OUT), .A1 (XNOR_1_1_NUM16_OUT), .A2 (XNOR_1_2_NUM16_OUT));

      wire XNOR_2_1_NUM16_OUT, XNOR_2_2_NUM16_OUT;
      NOR2_X1 XNOR_2_1_NUM16 (.ZN (XNOR_2_1_NUM16_OUT), .A1 (N80), .A2 (GND));
      NOR2_X1 XNOR_2_2_NUM16 (.ZN (XNOR_2_2_NUM16_OUT), .A1 (GND), .A2 (XNOR_1_3_NUM16_OUT));
      NOR2_X1 XNOR_2_3_NUM16 (.ZN (N295), .A1 (XNOR_2_1_NUM16_OUT), .A2 (XNOR_2_2_NUM16_OUT));
      wire XNOR_1_1_NUM17_OUT, XNOR_1_2_NUM17_OUT, XNOR_1_3_NUM17_OUT;
      NOR2_X1 XNOR_1_1_NUM17 (.ZN (XNOR_1_1_NUM17_OUT), .A1 (N59), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM17 (.ZN (XNOR_1_2_NUM17_OUT), .A1 (GND), .A2 (N36));
      NOR2_X1 XNOR_1_3_NUM17 (.ZN (XNOR_1_3_NUM17_OUT), .A1 (XNOR_1_1_NUM17_OUT), .A2 (XNOR_1_2_NUM17_OUT));

      wire XNOR_2_1_NUM17_OUT, XNOR_2_2_NUM17_OUT;
      NOR2_X1 XNOR_2_1_NUM17 (.ZN (XNOR_2_1_NUM17_OUT), .A1 (N42), .A2 (GND));
      NOR2_X1 XNOR_2_2_NUM17 (.ZN (XNOR_2_2_NUM17_OUT), .A1 (GND), .A2 (XNOR_1_3_NUM17_OUT));
      NOR2_X1 XNOR_2_3_NUM17 (.ZN (N296), .A1 (XNOR_2_1_NUM17_OUT), .A2 (XNOR_2_2_NUM17_OUT));
      wire XNOR_1_1_NUM18_OUT, XNOR_1_2_NUM18_OUT;
      NOR2_X1 XNOR_1_1_NUM18 (.ZN (XNOR_1_1_NUM18_OUT), .A1 (N85), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM18 (.ZN (XNOR_1_2_NUM18_OUT), .A1 (GND), .A2 (N86));
      NOR2_X1 XNOR_1_3_NUM18 (.ZN (N297), .A1 (XNOR_1_1_NUM18_OUT), .A2 (XNOR_1_2_NUM18_OUT));
      wire XNOR_1_NUM19_OUT;
      NOR2_X1 XNOR_1_NUM19 (.ZN (XNOR_1_NUM19_OUT), .A1 (N87), .A2 (N88));
      NOR2_X1 XNOR_2_NUM19 (.ZN (N298), .A1 (XNOR_1_NUM19_OUT), .A2 (GND));
      wire XNOR_1_1_NUM20_OUT, XNOR_1_2_NUM20_OUT, XNOR_1_3_NUM20_OUT;
      NOR2_X1 XNOR_1_1_NUM20 (.ZN (XNOR_1_1_NUM20_OUT), .A1 (N91), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM20 (.ZN (XNOR_1_2_NUM20_OUT), .A1 (GND), .A2 (N96));
      NOR2_X1 XNOR_1_3_NUM20 (.ZN (XNOR_1_3_NUM20_OUT), .A1 (XNOR_1_1_NUM20_OUT), .A2 (XNOR_1_2_NUM20_OUT));
      NOR2_X1 XNOR_1_4_NUM20 (.ZN (N301), .A1 (XNOR_1_3_NUM20_OUT), .A2 (GND));
      wire XNOR_1_NUM21_OUT;
      NOR2_X1 XNOR_1_NUM21 (.ZN (XNOR_1_NUM21_OUT), .A1 (N91), .A2 (N96));
      NOR2_X1 XNOR_2_NUM21 (.ZN (N302), .A1 (XNOR_1_NUM21_OUT), .A2 (GND));
      wire XNOR_1_1_NUM22_OUT, XNOR_1_2_NUM22_OUT, XNOR_1_3_NUM22_OUT;
      NOR2_X1 XNOR_1_1_NUM22 (.ZN (XNOR_1_1_NUM22_OUT), .A1 (N101), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM22 (.ZN (XNOR_1_2_NUM22_OUT), .A1 (GND), .A2 (N106));
      NOR2_X1 XNOR_1_3_NUM22 (.ZN (XNOR_1_3_NUM22_OUT), .A1 (XNOR_1_1_NUM22_OUT), .A2 (XNOR_1_2_NUM22_OUT));
      NOR2_X1 XNOR_1_4_NUM22 (.ZN (N303), .A1 (XNOR_1_3_NUM22_OUT), .A2 (GND));
      wire XNOR_1_NUM23_OUT;
      NOR2_X1 XNOR_1_NUM23 (.ZN (XNOR_1_NUM23_OUT), .A1 (N101), .A2 (N106));
      NOR2_X1 XNOR_2_NUM23 (.ZN (N304), .A1 (XNOR_1_NUM23_OUT), .A2 (GND));
      wire XNOR_1_1_NUM24_OUT, XNOR_1_2_NUM24_OUT, XNOR_1_3_NUM24_OUT;
      NOR2_X1 XNOR_1_1_NUM24 (.ZN (XNOR_1_1_NUM24_OUT), .A1 (N111), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM24 (.ZN (XNOR_1_2_NUM24_OUT), .A1 (GND), .A2 (N116));
      NOR2_X1 XNOR_1_3_NUM24 (.ZN (XNOR_1_3_NUM24_OUT), .A1 (XNOR_1_1_NUM24_OUT), .A2 (XNOR_1_2_NUM24_OUT));
      NOR2_X1 XNOR_1_4_NUM24 (.ZN (N305), .A1 (XNOR_1_3_NUM24_OUT), .A2 (GND));
      wire XNOR_1_NUM25_OUT;
      NOR2_X1 XNOR_1_NUM25 (.ZN (XNOR_1_NUM25_OUT), .A1 (N111), .A2 (N116));
      NOR2_X1 XNOR_2_NUM25 (.ZN (N306), .A1 (XNOR_1_NUM25_OUT), .A2 (GND));
      wire XNOR_1_1_NUM26_OUT, XNOR_1_2_NUM26_OUT, XNOR_1_3_NUM26_OUT;
      NOR2_X1 XNOR_1_1_NUM26 (.ZN (XNOR_1_1_NUM26_OUT), .A1 (N121), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM26 (.ZN (XNOR_1_2_NUM26_OUT), .A1 (GND), .A2 (N126));
      NOR2_X1 XNOR_1_3_NUM26 (.ZN (XNOR_1_3_NUM26_OUT), .A1 (XNOR_1_1_NUM26_OUT), .A2 (XNOR_1_2_NUM26_OUT));
      NOR2_X1 XNOR_1_4_NUM26 (.ZN (N307), .A1 (XNOR_1_3_NUM26_OUT), .A2 (GND));
      wire XNOR_1_NUM27_OUT;
      NOR2_X1 XNOR_1_NUM27 (.ZN (XNOR_1_NUM27_OUT), .A1 (N121), .A2 (N126));
      NOR2_X1 XNOR_2_NUM27 (.ZN (N308), .A1 (XNOR_1_NUM27_OUT), .A2 (GND));
      wire XNOR_1_1_NUM28_OUT, XNOR_1_2_NUM28_OUT;
      NOR2_X1 XNOR_1_1_NUM28 (.ZN (XNOR_1_1_NUM28_OUT), .A1 (N8), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM28 (.ZN (XNOR_1_2_NUM28_OUT), .A1 (GND), .A2 (N138));
      NOR2_X1 XNOR_1_3_NUM28 (.ZN (N309), .A1 (XNOR_1_1_NUM28_OUT), .A2 (XNOR_1_2_NUM28_OUT));
      NOR2_X1 XNOR_NUM29 (.ZN (N310), .A1 (N268), .A2 (GND));
      wire XNOR_1_1_NUM30_OUT, XNOR_1_2_NUM30_OUT;
      NOR2_X1 XNOR_1_1_NUM30 (.ZN (XNOR_1_1_NUM30_OUT), .A1 (N51), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM30 (.ZN (XNOR_1_2_NUM30_OUT), .A1 (GND), .A2 (N138));
      NOR2_X1 XNOR_1_3_NUM30 (.ZN (N316), .A1 (XNOR_1_1_NUM30_OUT), .A2 (XNOR_1_2_NUM30_OUT));
      wire XNOR_1_1_NUM31_OUT, XNOR_1_2_NUM31_OUT;
      NOR2_X1 XNOR_1_1_NUM31 (.ZN (XNOR_1_1_NUM31_OUT), .A1 (N17), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM31 (.ZN (XNOR_1_2_NUM31_OUT), .A1 (GND), .A2 (N138));
      NOR2_X1 XNOR_1_3_NUM31 (.ZN (N317), .A1 (XNOR_1_1_NUM31_OUT), .A2 (XNOR_1_2_NUM31_OUT));
      wire XNOR_1_1_NUM32_OUT, XNOR_1_2_NUM32_OUT;
      NOR2_X1 XNOR_1_1_NUM32 (.ZN (XNOR_1_1_NUM32_OUT), .A1 (N152), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM32 (.ZN (XNOR_1_2_NUM32_OUT), .A1 (GND), .A2 (N138));
      NOR2_X1 XNOR_1_3_NUM32 (.ZN (N318), .A1 (XNOR_1_1_NUM32_OUT), .A2 (XNOR_1_2_NUM32_OUT));
      wire XNOR_1_1_NUM33_OUT, XNOR_1_2_NUM33_OUT, XNOR_1_3_NUM33_OUT;
      NOR2_X1 XNOR_1_1_NUM33 (.ZN (XNOR_1_1_NUM33_OUT), .A1 (N59), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM33 (.ZN (XNOR_1_2_NUM33_OUT), .A1 (GND), .A2 (N156));
      NOR2_X1 XNOR_1_3_NUM33 (.ZN (XNOR_1_3_NUM33_OUT), .A1 (XNOR_1_1_NUM33_OUT), .A2 (XNOR_1_2_NUM33_OUT));
      NOR2_X1 XNOR_1_4_NUM33 (.ZN (N319), .A1 (XNOR_1_3_NUM33_OUT), .A2 (GND));
      NOR2_X1 XNOR_NUM34 (.ZN (N322), .A1 (N17), .A2 (N42));
      wire XNOR_1_1_NUM35_OUT, XNOR_1_2_NUM35_OUT;
      NOR2_X1 XNOR_1_1_NUM35 (.ZN (XNOR_1_1_NUM35_OUT), .A1 (N17), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM35 (.ZN (XNOR_1_2_NUM35_OUT), .A1 (GND), .A2 (N42));
      NOR2_X1 XNOR_1_3_NUM35 (.ZN (N323), .A1 (XNOR_1_1_NUM35_OUT), .A2 (XNOR_1_2_NUM35_OUT));
      wire XNOR_1_1_NUM36_OUT, XNOR_1_2_NUM36_OUT, XNOR_1_3_NUM36_OUT;
      NOR2_X1 XNOR_1_1_NUM36 (.ZN (XNOR_1_1_NUM36_OUT), .A1 (N159), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM36 (.ZN (XNOR_1_2_NUM36_OUT), .A1 (GND), .A2 (N165));
      NOR2_X1 XNOR_1_3_NUM36 (.ZN (XNOR_1_3_NUM36_OUT), .A1 (XNOR_1_1_NUM36_OUT), .A2 (XNOR_1_2_NUM36_OUT));
      NOR2_X1 XNOR_1_4_NUM36 (.ZN (N324), .A1 (XNOR_1_3_NUM36_OUT), .A2 (GND));
      wire XNOR_1_NUM37_OUT;
      NOR2_X1 XNOR_1_NUM37 (.ZN (XNOR_1_NUM37_OUT), .A1 (N159), .A2 (N165));
      NOR2_X1 XNOR_2_NUM37 (.ZN (N325), .A1 (XNOR_1_NUM37_OUT), .A2 (GND));
      wire XNOR_1_1_NUM38_OUT, XNOR_1_2_NUM38_OUT, XNOR_1_3_NUM38_OUT;
      NOR2_X1 XNOR_1_1_NUM38 (.ZN (XNOR_1_1_NUM38_OUT), .A1 (N171), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM38 (.ZN (XNOR_1_2_NUM38_OUT), .A1 (GND), .A2 (N177));
      NOR2_X1 XNOR_1_3_NUM38 (.ZN (XNOR_1_3_NUM38_OUT), .A1 (XNOR_1_1_NUM38_OUT), .A2 (XNOR_1_2_NUM38_OUT));
      NOR2_X1 XNOR_1_4_NUM38 (.ZN (N326), .A1 (XNOR_1_3_NUM38_OUT), .A2 (GND));
      wire XNOR_1_NUM39_OUT;
      NOR2_X1 XNOR_1_NUM39 (.ZN (XNOR_1_NUM39_OUT), .A1 (N171), .A2 (N177));
      NOR2_X1 XNOR_2_NUM39 (.ZN (N327), .A1 (XNOR_1_NUM39_OUT), .A2 (GND));
      wire XNOR_1_1_NUM40_OUT, XNOR_1_2_NUM40_OUT, XNOR_1_3_NUM40_OUT;
      NOR2_X1 XNOR_1_1_NUM40 (.ZN (XNOR_1_1_NUM40_OUT), .A1 (N183), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM40 (.ZN (XNOR_1_2_NUM40_OUT), .A1 (GND), .A2 (N189));
      NOR2_X1 XNOR_1_3_NUM40 (.ZN (XNOR_1_3_NUM40_OUT), .A1 (XNOR_1_1_NUM40_OUT), .A2 (XNOR_1_2_NUM40_OUT));
      NOR2_X1 XNOR_1_4_NUM40 (.ZN (N328), .A1 (XNOR_1_3_NUM40_OUT), .A2 (GND));
      wire XNOR_1_NUM41_OUT;
      NOR2_X1 XNOR_1_NUM41 (.ZN (XNOR_1_NUM41_OUT), .A1 (N183), .A2 (N189));
      NOR2_X1 XNOR_2_NUM41 (.ZN (N329), .A1 (XNOR_1_NUM41_OUT), .A2 (GND));
      wire XNOR_1_1_NUM42_OUT, XNOR_1_2_NUM42_OUT, XNOR_1_3_NUM42_OUT;
      NOR2_X1 XNOR_1_1_NUM42 (.ZN (XNOR_1_1_NUM42_OUT), .A1 (N195), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM42 (.ZN (XNOR_1_2_NUM42_OUT), .A1 (GND), .A2 (N201));
      NOR2_X1 XNOR_1_3_NUM42 (.ZN (XNOR_1_3_NUM42_OUT), .A1 (XNOR_1_1_NUM42_OUT), .A2 (XNOR_1_2_NUM42_OUT));
      NOR2_X1 XNOR_1_4_NUM42 (.ZN (N330), .A1 (XNOR_1_3_NUM42_OUT), .A2 (GND));
      wire XNOR_1_NUM43_OUT;
      NOR2_X1 XNOR_1_NUM43 (.ZN (XNOR_1_NUM43_OUT), .A1 (N195), .A2 (N201));
      NOR2_X1 XNOR_2_NUM43 (.ZN (N331), .A1 (XNOR_1_NUM43_OUT), .A2 (GND));
      wire XNOR_1_1_NUM44_OUT, XNOR_1_2_NUM44_OUT;
      NOR2_X1 XNOR_1_1_NUM44 (.ZN (XNOR_1_1_NUM44_OUT), .A1 (N210), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM44 (.ZN (XNOR_1_2_NUM44_OUT), .A1 (GND), .A2 (N91));
      NOR2_X1 XNOR_1_3_NUM44 (.ZN (N332), .A1 (XNOR_1_1_NUM44_OUT), .A2 (XNOR_1_2_NUM44_OUT));
      wire XNOR_1_1_NUM45_OUT, XNOR_1_2_NUM45_OUT;
      NOR2_X1 XNOR_1_1_NUM45 (.ZN (XNOR_1_1_NUM45_OUT), .A1 (N210), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM45 (.ZN (XNOR_1_2_NUM45_OUT), .A1 (GND), .A2 (N96));
      NOR2_X1 XNOR_1_3_NUM45 (.ZN (N333), .A1 (XNOR_1_1_NUM45_OUT), .A2 (XNOR_1_2_NUM45_OUT));
      wire XNOR_1_1_NUM46_OUT, XNOR_1_2_NUM46_OUT;
      NOR2_X1 XNOR_1_1_NUM46 (.ZN (XNOR_1_1_NUM46_OUT), .A1 (N210), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM46 (.ZN (XNOR_1_2_NUM46_OUT), .A1 (GND), .A2 (N101));
      NOR2_X1 XNOR_1_3_NUM46 (.ZN (N334), .A1 (XNOR_1_1_NUM46_OUT), .A2 (XNOR_1_2_NUM46_OUT));
      wire XNOR_1_1_NUM47_OUT, XNOR_1_2_NUM47_OUT;
      NOR2_X1 XNOR_1_1_NUM47 (.ZN (XNOR_1_1_NUM47_OUT), .A1 (N210), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM47 (.ZN (XNOR_1_2_NUM47_OUT), .A1 (GND), .A2 (N106));
      NOR2_X1 XNOR_1_3_NUM47 (.ZN (N335), .A1 (XNOR_1_1_NUM47_OUT), .A2 (XNOR_1_2_NUM47_OUT));
      wire XNOR_1_1_NUM48_OUT, XNOR_1_2_NUM48_OUT;
      NOR2_X1 XNOR_1_1_NUM48 (.ZN (XNOR_1_1_NUM48_OUT), .A1 (N210), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM48 (.ZN (XNOR_1_2_NUM48_OUT), .A1 (GND), .A2 (N111));
      NOR2_X1 XNOR_1_3_NUM48 (.ZN (N336), .A1 (XNOR_1_1_NUM48_OUT), .A2 (XNOR_1_2_NUM48_OUT));
      wire XNOR_1_1_NUM49_OUT, XNOR_1_2_NUM49_OUT;
      NOR2_X1 XNOR_1_1_NUM49 (.ZN (XNOR_1_1_NUM49_OUT), .A1 (N255), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM49 (.ZN (XNOR_1_2_NUM49_OUT), .A1 (GND), .A2 (N259));
      NOR2_X1 XNOR_1_3_NUM49 (.ZN (N337), .A1 (XNOR_1_1_NUM49_OUT), .A2 (XNOR_1_2_NUM49_OUT));
      wire XNOR_1_1_NUM50_OUT, XNOR_1_2_NUM50_OUT;
      NOR2_X1 XNOR_1_1_NUM50 (.ZN (XNOR_1_1_NUM50_OUT), .A1 (N210), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM50 (.ZN (XNOR_1_2_NUM50_OUT), .A1 (GND), .A2 (N116));
      NOR2_X1 XNOR_1_3_NUM50 (.ZN (N338), .A1 (XNOR_1_1_NUM50_OUT), .A2 (XNOR_1_2_NUM50_OUT));
      wire XNOR_1_1_NUM51_OUT, XNOR_1_2_NUM51_OUT;
      NOR2_X1 XNOR_1_1_NUM51 (.ZN (XNOR_1_1_NUM51_OUT), .A1 (N255), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM51 (.ZN (XNOR_1_2_NUM51_OUT), .A1 (GND), .A2 (N260));
      NOR2_X1 XNOR_1_3_NUM51 (.ZN (N339), .A1 (XNOR_1_1_NUM51_OUT), .A2 (XNOR_1_2_NUM51_OUT));
      wire XNOR_1_1_NUM52_OUT, XNOR_1_2_NUM52_OUT;
      NOR2_X1 XNOR_1_1_NUM52 (.ZN (XNOR_1_1_NUM52_OUT), .A1 (N210), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM52 (.ZN (XNOR_1_2_NUM52_OUT), .A1 (GND), .A2 (N121));
      NOR2_X1 XNOR_1_3_NUM52 (.ZN (N340), .A1 (XNOR_1_1_NUM52_OUT), .A2 (XNOR_1_2_NUM52_OUT));
      wire XNOR_1_1_NUM53_OUT, XNOR_1_2_NUM53_OUT;
      NOR2_X1 XNOR_1_1_NUM53 (.ZN (XNOR_1_1_NUM53_OUT), .A1 (N255), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM53 (.ZN (XNOR_1_2_NUM53_OUT), .A1 (GND), .A2 (N267));
      NOR2_X1 XNOR_1_3_NUM53 (.ZN (N341), .A1 (XNOR_1_1_NUM53_OUT), .A2 (XNOR_1_2_NUM53_OUT));
      NOR2_X1 XNOR_NUM54 (.ZN (N342), .A1 (N269), .A2 (GND));
      NOR2_X1 XNOR_NUM55 (.ZN (N343), .A1 (N273), .A2 (GND));
      wire XNOR_1_NUM56_OUT;
      NOR2_X1 XNOR_1_NUM56 (.ZN (XNOR_1_NUM56_OUT), .A1 (N270), .A2 (N273));
      NOR2_X1 XNOR_2_NUM56 (.ZN (N344), .A1 (XNOR_1_NUM56_OUT), .A2 (GND));
      NOR2_X1 XNOR_NUM57 (.ZN (N345), .A1 (N276), .A2 (GND));
      NOR2_X1 XNOR_NUM58 (.ZN (N346), .A1 (N276), .A2 (GND));
      NOR2_X1 XNOR_NUM59 (.ZN (N347), .A1 (N279), .A2 (GND));
      NOR2_X1 XNOR_NUM60 (.ZN (N348), .A1 (N280), .A2 (N284));
      wire XNOR_1_NUM61_OUT;
      NOR2_X1 XNOR_1_NUM61 (.ZN (XNOR_1_NUM61_OUT), .A1 (N280), .A2 (N285));
      NOR2_X1 XNOR_2_NUM61 (.ZN (N349), .A1 (XNOR_1_NUM61_OUT), .A2 (GND));
      wire XNOR_1_NUM62_OUT;
      NOR2_X1 XNOR_1_NUM62 (.ZN (XNOR_1_NUM62_OUT), .A1 (N280), .A2 (N286));
      NOR2_X1 XNOR_2_NUM62 (.ZN (N350), .A1 (XNOR_1_NUM62_OUT), .A2 (GND));
      NOR2_X1 XNOR_NUM63 (.ZN (N351), .A1 (N293), .A2 (GND));
      NOR2_X1 XNOR_NUM64 (.ZN (N352), .A1 (N294), .A2 (GND));
      NOR2_X1 XNOR_NUM65 (.ZN (N353), .A1 (N295), .A2 (GND));
      NOR2_X1 XNOR_NUM66 (.ZN (N354), .A1 (N296), .A2 (GND));
      wire XNOR_1_1_NUM67_OUT, XNOR_1_2_NUM67_OUT, XNOR_1_3_NUM67_OUT;
      NOR2_X1 XNOR_1_1_NUM67 (.ZN (XNOR_1_1_NUM67_OUT), .A1 (N89), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM67 (.ZN (XNOR_1_2_NUM67_OUT), .A1 (GND), .A2 (N298));
      NOR2_X1 XNOR_1_3_NUM67 (.ZN (XNOR_1_3_NUM67_OUT), .A1 (XNOR_1_1_NUM67_OUT), .A2 (XNOR_1_2_NUM67_OUT));
      NOR2_X1 XNOR_1_4_NUM67 (.ZN (N355), .A1 (XNOR_1_3_NUM67_OUT), .A2 (GND));
      wire XNOR_1_1_NUM68_OUT, XNOR_1_2_NUM68_OUT;
      NOR2_X1 XNOR_1_1_NUM68 (.ZN (XNOR_1_1_NUM68_OUT), .A1 (N90), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM68 (.ZN (XNOR_1_2_NUM68_OUT), .A1 (GND), .A2 (N298));
      NOR2_X1 XNOR_1_3_NUM68 (.ZN (N356), .A1 (XNOR_1_1_NUM68_OUT), .A2 (XNOR_1_2_NUM68_OUT));
      wire XNOR_1_1_NUM69_OUT, XNOR_1_2_NUM69_OUT, XNOR_1_3_NUM69_OUT;
      NOR2_X1 XNOR_1_1_NUM69 (.ZN (XNOR_1_1_NUM69_OUT), .A1 (N301), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM69 (.ZN (XNOR_1_2_NUM69_OUT), .A1 (GND), .A2 (N302));
      NOR2_X1 XNOR_1_3_NUM69 (.ZN (XNOR_1_3_NUM69_OUT), .A1 (XNOR_1_1_NUM69_OUT), .A2 (XNOR_1_2_NUM69_OUT));
      NOR2_X1 XNOR_1_4_NUM69 (.ZN (N357), .A1 (XNOR_1_3_NUM69_OUT), .A2 (GND));
      wire XNOR_1_1_NUM70_OUT, XNOR_1_2_NUM70_OUT, XNOR_1_3_NUM70_OUT;
      NOR2_X1 XNOR_1_1_NUM70 (.ZN (XNOR_1_1_NUM70_OUT), .A1 (N303), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM70 (.ZN (XNOR_1_2_NUM70_OUT), .A1 (GND), .A2 (N304));
      NOR2_X1 XNOR_1_3_NUM70 (.ZN (XNOR_1_3_NUM70_OUT), .A1 (XNOR_1_1_NUM70_OUT), .A2 (XNOR_1_2_NUM70_OUT));
      NOR2_X1 XNOR_1_4_NUM70 (.ZN (N360), .A1 (XNOR_1_3_NUM70_OUT), .A2 (GND));
      wire XNOR_1_1_NUM71_OUT, XNOR_1_2_NUM71_OUT, XNOR_1_3_NUM71_OUT;
      NOR2_X1 XNOR_1_1_NUM71 (.ZN (XNOR_1_1_NUM71_OUT), .A1 (N305), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM71 (.ZN (XNOR_1_2_NUM71_OUT), .A1 (GND), .A2 (N306));
      NOR2_X1 XNOR_1_3_NUM71 (.ZN (XNOR_1_3_NUM71_OUT), .A1 (XNOR_1_1_NUM71_OUT), .A2 (XNOR_1_2_NUM71_OUT));
      NOR2_X1 XNOR_1_4_NUM71 (.ZN (N363), .A1 (XNOR_1_3_NUM71_OUT), .A2 (GND));
      wire XNOR_1_1_NUM72_OUT, XNOR_1_2_NUM72_OUT, XNOR_1_3_NUM72_OUT;
      NOR2_X1 XNOR_1_1_NUM72 (.ZN (XNOR_1_1_NUM72_OUT), .A1 (N307), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM72 (.ZN (XNOR_1_2_NUM72_OUT), .A1 (GND), .A2 (N308));
      NOR2_X1 XNOR_1_3_NUM72 (.ZN (XNOR_1_3_NUM72_OUT), .A1 (XNOR_1_1_NUM72_OUT), .A2 (XNOR_1_2_NUM72_OUT));
      NOR2_X1 XNOR_1_4_NUM72 (.ZN (N366), .A1 (XNOR_1_3_NUM72_OUT), .A2 (GND));
      NOR2_X1 XNOR_NUM73 (.ZN (N369), .A1 (N310), .A2 (GND));
      NOR2_X1 XNOR_NUM74 (.ZN (N375), .A1 (N322), .A2 (N323));
      wire XNOR_1_1_NUM75_OUT, XNOR_1_2_NUM75_OUT, XNOR_1_3_NUM75_OUT;
      NOR2_X1 XNOR_1_1_NUM75 (.ZN (XNOR_1_1_NUM75_OUT), .A1 (N324), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM75 (.ZN (XNOR_1_2_NUM75_OUT), .A1 (GND), .A2 (N325));
      NOR2_X1 XNOR_1_3_NUM75 (.ZN (XNOR_1_3_NUM75_OUT), .A1 (XNOR_1_1_NUM75_OUT), .A2 (XNOR_1_2_NUM75_OUT));
      NOR2_X1 XNOR_1_4_NUM75 (.ZN (N376), .A1 (XNOR_1_3_NUM75_OUT), .A2 (GND));
      wire XNOR_1_1_NUM76_OUT, XNOR_1_2_NUM76_OUT, XNOR_1_3_NUM76_OUT;
      NOR2_X1 XNOR_1_1_NUM76 (.ZN (XNOR_1_1_NUM76_OUT), .A1 (N326), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM76 (.ZN (XNOR_1_2_NUM76_OUT), .A1 (GND), .A2 (N327));
      NOR2_X1 XNOR_1_3_NUM76 (.ZN (XNOR_1_3_NUM76_OUT), .A1 (XNOR_1_1_NUM76_OUT), .A2 (XNOR_1_2_NUM76_OUT));
      NOR2_X1 XNOR_1_4_NUM76 (.ZN (N379), .A1 (XNOR_1_3_NUM76_OUT), .A2 (GND));
      wire XNOR_1_1_NUM77_OUT, XNOR_1_2_NUM77_OUT, XNOR_1_3_NUM77_OUT;
      NOR2_X1 XNOR_1_1_NUM77 (.ZN (XNOR_1_1_NUM77_OUT), .A1 (N328), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM77 (.ZN (XNOR_1_2_NUM77_OUT), .A1 (GND), .A2 (N329));
      NOR2_X1 XNOR_1_3_NUM77 (.ZN (XNOR_1_3_NUM77_OUT), .A1 (XNOR_1_1_NUM77_OUT), .A2 (XNOR_1_2_NUM77_OUT));
      NOR2_X1 XNOR_1_4_NUM77 (.ZN (N382), .A1 (XNOR_1_3_NUM77_OUT), .A2 (GND));
      wire XNOR_1_1_NUM78_OUT, XNOR_1_2_NUM78_OUT, XNOR_1_3_NUM78_OUT;
      NOR2_X1 XNOR_1_1_NUM78 (.ZN (XNOR_1_1_NUM78_OUT), .A1 (N330), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM78 (.ZN (XNOR_1_2_NUM78_OUT), .A1 (GND), .A2 (N331));
      NOR2_X1 XNOR_1_3_NUM78 (.ZN (XNOR_1_3_NUM78_OUT), .A1 (XNOR_1_1_NUM78_OUT), .A2 (XNOR_1_2_NUM78_OUT));
      NOR2_X1 XNOR_1_4_NUM78 (.ZN (N385), .A1 (XNOR_1_3_NUM78_OUT), .A2 (GND));
      wire XNOR_1_1_NUM79_OUT;
      NOR2_X1 XNOR_1_1_NUM79 (.ZN (XNOR_1_1_NUM79_OUT), .A1 (N290), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM79 (.ZN (N388), .A1 (XNOR_1_1_NUM79_OUT), .A2 (GND));
      wire XNOR_1_1_NUM80_OUT;
      NOR2_X1 XNOR_1_1_NUM80 (.ZN (XNOR_1_1_NUM80_OUT), .A1 (N291), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM80 (.ZN (N389), .A1 (XNOR_1_1_NUM80_OUT), .A2 (GND));
      wire XNOR_1_1_NUM81_OUT;
      NOR2_X1 XNOR_1_1_NUM81 (.ZN (XNOR_1_1_NUM81_OUT), .A1 (N292), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM81 (.ZN (N390), .A1 (XNOR_1_1_NUM81_OUT), .A2 (GND));
      wire XNOR_1_1_NUM82_OUT;
      NOR2_X1 XNOR_1_1_NUM82 (.ZN (XNOR_1_1_NUM82_OUT), .A1 (N297), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM82 (.ZN (N391), .A1 (XNOR_1_1_NUM82_OUT), .A2 (GND));
      wire XNOR_1_NUM83_OUT;
      NOR2_X1 XNOR_1_NUM83 (.ZN (XNOR_1_NUM83_OUT), .A1 (N270), .A2 (N343));
      NOR2_X1 XNOR_2_NUM83 (.ZN (N392), .A1 (XNOR_1_NUM83_OUT), .A2 (GND));
      NOR2_X1 XNOR_NUM84 (.ZN (N393), .A1 (N345), .A2 (GND));
      NOR2_X1 XNOR_NUM85 (.ZN (N399), .A1 (N346), .A2 (GND));
      wire XNOR_1_1_NUM86_OUT, XNOR_1_2_NUM86_OUT;
      NOR2_X1 XNOR_1_1_NUM86 (.ZN (XNOR_1_1_NUM86_OUT), .A1 (N348), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM86 (.ZN (XNOR_1_2_NUM86_OUT), .A1 (GND), .A2 (N73));
      NOR2_X1 XNOR_1_3_NUM86 (.ZN (N400), .A1 (XNOR_1_1_NUM86_OUT), .A2 (XNOR_1_2_NUM86_OUT));
      NOR2_X1 XNOR_NUM87 (.ZN (N401), .A1 (N349), .A2 (GND));
      NOR2_X1 XNOR_NUM88 (.ZN (N402), .A1 (N350), .A2 (GND));
      NOR2_X1 XNOR_NUM89 (.ZN (N403), .A1 (N355), .A2 (GND));
      NOR2_X1 XNOR_NUM90 (.ZN (N404), .A1 (N357), .A2 (GND));
      NOR2_X1 XNOR_NUM91 (.ZN (N405), .A1 (N360), .A2 (GND));
      wire XNOR_1_1_NUM92_OUT, XNOR_1_2_NUM92_OUT;
      NOR2_X1 XNOR_1_1_NUM92 (.ZN (XNOR_1_1_NUM92_OUT), .A1 (N357), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM92 (.ZN (XNOR_1_2_NUM92_OUT), .A1 (GND), .A2 (N360));
      NOR2_X1 XNOR_1_3_NUM92 (.ZN (N406), .A1 (XNOR_1_1_NUM92_OUT), .A2 (XNOR_1_2_NUM92_OUT));
      NOR2_X1 XNOR_NUM93 (.ZN (N407), .A1 (N363), .A2 (GND));
      NOR2_X1 XNOR_NUM94 (.ZN (N408), .A1 (N366), .A2 (GND));
      wire XNOR_1_1_NUM95_OUT, XNOR_1_2_NUM95_OUT;
      NOR2_X1 XNOR_1_1_NUM95 (.ZN (XNOR_1_1_NUM95_OUT), .A1 (N363), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM95 (.ZN (XNOR_1_2_NUM95_OUT), .A1 (GND), .A2 (N366));
      NOR2_X1 XNOR_1_3_NUM95 (.ZN (N409), .A1 (XNOR_1_1_NUM95_OUT), .A2 (XNOR_1_2_NUM95_OUT));
      wire XNOR_1_1_NUM96_OUT, XNOR_1_2_NUM96_OUT, XNOR_1_3_NUM96_OUT;
      NOR2_X1 XNOR_1_1_NUM96 (.ZN (XNOR_1_1_NUM96_OUT), .A1 (N347), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM96 (.ZN (XNOR_1_2_NUM96_OUT), .A1 (GND), .A2 (N352));
      NOR2_X1 XNOR_1_3_NUM96 (.ZN (XNOR_1_3_NUM96_OUT), .A1 (XNOR_1_1_NUM96_OUT), .A2 (XNOR_1_2_NUM96_OUT));
      NOR2_X1 XNOR_1_4_NUM96 (.ZN (N410), .A1 (XNOR_1_3_NUM96_OUT), .A2 (GND));
      NOR2_X1 XNOR_NUM97 (.ZN (N411), .A1 (N376), .A2 (GND));
      NOR2_X1 XNOR_NUM98 (.ZN (N412), .A1 (N379), .A2 (GND));
      wire XNOR_1_1_NUM99_OUT, XNOR_1_2_NUM99_OUT;
      NOR2_X1 XNOR_1_1_NUM99 (.ZN (XNOR_1_1_NUM99_OUT), .A1 (N376), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM99 (.ZN (XNOR_1_2_NUM99_OUT), .A1 (GND), .A2 (N379));
      NOR2_X1 XNOR_1_3_NUM99 (.ZN (N413), .A1 (XNOR_1_1_NUM99_OUT), .A2 (XNOR_1_2_NUM99_OUT));
      NOR2_X1 XNOR_NUM100 (.ZN (N414), .A1 (N382), .A2 (GND));
      NOR2_X1 XNOR_NUM101 (.ZN (N415), .A1 (N385), .A2 (GND));
      wire XNOR_1_1_NUM102_OUT, XNOR_1_2_NUM102_OUT;
      NOR2_X1 XNOR_1_1_NUM102 (.ZN (XNOR_1_1_NUM102_OUT), .A1 (N382), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM102 (.ZN (XNOR_1_2_NUM102_OUT), .A1 (GND), .A2 (N385));
      NOR2_X1 XNOR_1_3_NUM102 (.ZN (N416), .A1 (XNOR_1_1_NUM102_OUT), .A2 (XNOR_1_2_NUM102_OUT));
      wire XNOR_1_1_NUM103_OUT, XNOR_1_2_NUM103_OUT;
      NOR2_X1 XNOR_1_1_NUM103 (.ZN (XNOR_1_1_NUM103_OUT), .A1 (N210), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM103 (.ZN (XNOR_1_2_NUM103_OUT), .A1 (GND), .A2 (N369));
      NOR2_X1 XNOR_1_3_NUM103 (.ZN (N417), .A1 (XNOR_1_1_NUM103_OUT), .A2 (XNOR_1_2_NUM103_OUT));
      wire XNOR_1_1_NUM104_OUT;
      NOR2_X1 XNOR_1_1_NUM104 (.ZN (XNOR_1_1_NUM104_OUT), .A1 (N342), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM104 (.ZN (N418), .A1 (XNOR_1_1_NUM104_OUT), .A2 (GND));
      wire XNOR_1_1_NUM105_OUT;
      NOR2_X1 XNOR_1_1_NUM105 (.ZN (XNOR_1_1_NUM105_OUT), .A1 (N344), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM105 (.ZN (N419), .A1 (XNOR_1_1_NUM105_OUT), .A2 (GND));
      wire XNOR_1_1_NUM106_OUT;
      NOR2_X1 XNOR_1_1_NUM106 (.ZN (XNOR_1_1_NUM106_OUT), .A1 (N351), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM106 (.ZN (N420), .A1 (XNOR_1_1_NUM106_OUT), .A2 (GND));
      wire XNOR_1_1_NUM107_OUT;
      NOR2_X1 XNOR_1_1_NUM107 (.ZN (XNOR_1_1_NUM107_OUT), .A1 (N353), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM107 (.ZN (N421), .A1 (XNOR_1_1_NUM107_OUT), .A2 (GND));
      wire XNOR_1_1_NUM108_OUT;
      NOR2_X1 XNOR_1_1_NUM108 (.ZN (XNOR_1_1_NUM108_OUT), .A1 (N354), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM108 (.ZN (N422), .A1 (XNOR_1_1_NUM108_OUT), .A2 (GND));
      wire XNOR_1_1_NUM109_OUT;
      NOR2_X1 XNOR_1_1_NUM109 (.ZN (XNOR_1_1_NUM109_OUT), .A1 (N356), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM109 (.ZN (N423), .A1 (XNOR_1_1_NUM109_OUT), .A2 (GND));
      NOR2_X1 XNOR_NUM110 (.ZN (N424), .A1 (N400), .A2 (GND));
      wire XNOR_1_1_NUM111_OUT, XNOR_1_2_NUM111_OUT;
      NOR2_X1 XNOR_1_1_NUM111 (.ZN (XNOR_1_1_NUM111_OUT), .A1 (N404), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM111 (.ZN (XNOR_1_2_NUM111_OUT), .A1 (GND), .A2 (N405));
      NOR2_X1 XNOR_1_3_NUM111 (.ZN (N425), .A1 (XNOR_1_1_NUM111_OUT), .A2 (XNOR_1_2_NUM111_OUT));
      wire XNOR_1_1_NUM112_OUT, XNOR_1_2_NUM112_OUT;
      NOR2_X1 XNOR_1_1_NUM112 (.ZN (XNOR_1_1_NUM112_OUT), .A1 (N407), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM112 (.ZN (XNOR_1_2_NUM112_OUT), .A1 (GND), .A2 (N408));
      NOR2_X1 XNOR_1_3_NUM112 (.ZN (N426), .A1 (XNOR_1_1_NUM112_OUT), .A2 (XNOR_1_2_NUM112_OUT));
      wire XNOR_1_1_NUM113_OUT, XNOR_1_2_NUM113_OUT, XNOR_1_3_NUM113_OUT;
      NOR2_X1 XNOR_1_1_NUM113 (.ZN (XNOR_1_1_NUM113_OUT), .A1 (N319), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM113 (.ZN (XNOR_1_2_NUM113_OUT), .A1 (GND), .A2 (N393));
      NOR2_X1 XNOR_1_3_NUM113 (.ZN (XNOR_1_3_NUM113_OUT), .A1 (XNOR_1_1_NUM113_OUT), .A2 (XNOR_1_2_NUM113_OUT));

      wire XNOR_2_1_NUM113_OUT, XNOR_2_2_NUM113_OUT;
      NOR2_X1 XNOR_2_1_NUM113 (.ZN (XNOR_2_1_NUM113_OUT), .A1 (N55), .A2 (GND));
      NOR2_X1 XNOR_2_2_NUM113 (.ZN (XNOR_2_2_NUM113_OUT), .A1 (GND), .A2 (XNOR_1_3_NUM113_OUT));
      NOR2_X1 XNOR_2_3_NUM113 (.ZN (N427), .A1 (XNOR_2_1_NUM113_OUT), .A2 (XNOR_2_2_NUM113_OUT));
      wire XNOR_1_1_NUM114_OUT, XNOR_1_2_NUM114_OUT, XNOR_1_3_NUM114_OUT;
      NOR2_X1 XNOR_1_1_NUM114 (.ZN (XNOR_1_1_NUM114_OUT), .A1 (N393), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM114 (.ZN (XNOR_1_2_NUM114_OUT), .A1 (GND), .A2 (N17));
      NOR2_X1 XNOR_1_3_NUM114 (.ZN (XNOR_1_3_NUM114_OUT), .A1 (XNOR_1_1_NUM114_OUT), .A2 (XNOR_1_2_NUM114_OUT));

      wire XNOR_2_1_NUM114_OUT, XNOR_2_2_NUM114_OUT;
      NOR2_X1 XNOR_2_1_NUM114 (.ZN (XNOR_2_1_NUM114_OUT), .A1 (N287), .A2 (GND));
      NOR2_X1 XNOR_2_2_NUM114 (.ZN (XNOR_2_2_NUM114_OUT), .A1 (GND), .A2 (XNOR_1_3_NUM114_OUT));
      NOR2_X1 XNOR_2_3_NUM114 (.ZN (N432), .A1 (XNOR_2_1_NUM114_OUT), .A2 (XNOR_2_2_NUM114_OUT));
      wire XNOR_1_1_NUM115_OUT, XNOR_1_2_NUM115_OUT, XNOR_1_3_NUM115_OUT;
      NOR2_X1 XNOR_1_1_NUM115 (.ZN (XNOR_1_1_NUM115_OUT), .A1 (N393), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM115 (.ZN (XNOR_1_2_NUM115_OUT), .A1 (GND), .A2 (N287));
      NOR2_X1 XNOR_1_3_NUM115 (.ZN (XNOR_1_3_NUM115_OUT), .A1 (XNOR_1_1_NUM115_OUT), .A2 (XNOR_1_2_NUM115_OUT));

      wire XNOR_2_1_NUM115_OUT, XNOR_2_2_NUM115_OUT, XNOR_2_3_NUM115_OUT;
      NOR2_X1 XNOR_2_1_NUM115 (.ZN (XNOR_2_1_NUM115_OUT), .A1 (N55), .A2 (GND));
      NOR2_X1 XNOR_2_2_NUM115 (.ZN (XNOR_2_2_NUM115_OUT), .A1 (GND), .A2 (XNOR_1_3_NUM115_OUT));
      NOR2_X1 XNOR_2_3_NUM115 (.ZN (XNOR_2_3_NUM115_OUT), .A1 (XNOR_2_1_NUM115_OUT), .A2 (XNOR_2_2_NUM115_OUT));

      NOR2_X1 XNOR_3_1_NUM115 (.ZN (N437), .A1 (XNOR_2_3_NUM115_OUT), .A2 (GND));
      wire XNOR_1_1_NUM116_OUT, XNOR_1_2_NUM116_OUT, XNOR_1_3_NUM116_OUT;
      NOR2_X1 XNOR_1_1_NUM116 (.ZN (XNOR_1_1_NUM116_OUT), .A1 (N375), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM116 (.ZN (XNOR_1_2_NUM116_OUT), .A1 (GND), .A2 (N59));
      NOR2_X1 XNOR_1_3_NUM116 (.ZN (XNOR_1_3_NUM116_OUT), .A1 (XNOR_1_1_NUM116_OUT), .A2 (XNOR_1_2_NUM116_OUT));

      wire XNOR_2_1_NUM116_OUT, XNOR_2_2_NUM116_OUT, XNOR_2_3_NUM116_OUT;
      NOR2_X1 XNOR_2_1_NUM116 (.ZN (XNOR_2_1_NUM116_OUT), .A1 (N156), .A2 (GND));
      NOR2_X1 XNOR_2_2_NUM116 (.ZN (XNOR_2_2_NUM116_OUT), .A1 (GND), .A2 (N393));
      NOR2_X1 XNOR_2_3_NUM116 (.ZN (XNOR_2_3_NUM116_OUT), .A1 (XNOR_2_1_NUM116_OUT), .A2 (XNOR_2_2_NUM116_OUT));

      wire XNOR_3_1_NUM116_OUT, XNOR_3_2_NUM116_OUT, XNOR_3_3_NUM116_OUT;
      NOR2_X1 XNOR_3_1_NUM116 (.ZN (XNOR_3_1_NUM116_OUT), .A1 (XNOR_1_3_NUM116_OUT), .A2 (GND));
      NOR2_X1 XNOR_3_2_NUM116 (.ZN (XNOR_3_2_NUM116_OUT), .A1 (GND), .A2 (XNOR_2_3_NUM116_OUT));
      NOR2_X1 XNOR_3_3_NUM116 (.ZN (XNOR_3_3_NUM116_OUT), .A1 (XNOR_3_1_NUM116_OUT), .A2 (XNOR_3_2_NUM116_OUT));

      NOR2_X1 XNOR_4_1_NUM116 (.ZN (N442), .A1 (XNOR_3_3_NUM116_OUT), .A2 (GND));
      wire XNOR_1_1_NUM117_OUT, XNOR_1_2_NUM117_OUT, XNOR_1_3_NUM117_OUT;
      NOR2_X1 XNOR_1_1_NUM117 (.ZN (XNOR_1_1_NUM117_OUT), .A1 (N393), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM117 (.ZN (XNOR_1_2_NUM117_OUT), .A1 (GND), .A2 (N319));
      NOR2_X1 XNOR_1_3_NUM117 (.ZN (XNOR_1_3_NUM117_OUT), .A1 (XNOR_1_1_NUM117_OUT), .A2 (XNOR_1_2_NUM117_OUT));

      wire XNOR_2_1_NUM117_OUT, XNOR_2_2_NUM117_OUT, XNOR_2_3_NUM117_OUT;
      NOR2_X1 XNOR_2_1_NUM117 (.ZN (XNOR_2_1_NUM117_OUT), .A1 (N17), .A2 (GND));
      NOR2_X1 XNOR_2_2_NUM117 (.ZN (XNOR_2_2_NUM117_OUT), .A1 (GND), .A2 (XNOR_1_3_NUM117_OUT));
      NOR2_X1 XNOR_2_3_NUM117 (.ZN (XNOR_2_3_NUM117_OUT), .A1 (XNOR_2_1_NUM117_OUT), .A2 (XNOR_2_2_NUM117_OUT));

      NOR2_X1 XNOR_3_1_NUM117 (.ZN (N443), .A1 (XNOR_2_3_NUM117_OUT), .A2 (GND));
      wire XNOR_1_1_NUM118_OUT, XNOR_1_2_NUM118_OUT;
      NOR2_X1 XNOR_1_1_NUM118 (.ZN (XNOR_1_1_NUM118_OUT), .A1 (N411), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM118 (.ZN (XNOR_1_2_NUM118_OUT), .A1 (GND), .A2 (N412));
      NOR2_X1 XNOR_1_3_NUM118 (.ZN (N444), .A1 (XNOR_1_1_NUM118_OUT), .A2 (XNOR_1_2_NUM118_OUT));
      wire XNOR_1_1_NUM119_OUT, XNOR_1_2_NUM119_OUT;
      NOR2_X1 XNOR_1_1_NUM119 (.ZN (XNOR_1_1_NUM119_OUT), .A1 (N414), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM119 (.ZN (XNOR_1_2_NUM119_OUT), .A1 (GND), .A2 (N415));
      NOR2_X1 XNOR_1_3_NUM119 (.ZN (N445), .A1 (XNOR_1_1_NUM119_OUT), .A2 (XNOR_1_2_NUM119_OUT));
      wire XNOR_1_1_NUM120_OUT;
      NOR2_X1 XNOR_1_1_NUM120 (.ZN (XNOR_1_1_NUM120_OUT), .A1 (N392), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM120 (.ZN (N446), .A1 (XNOR_1_1_NUM120_OUT), .A2 (GND));
      wire XNOR_1_1_NUM121_OUT;
      NOR2_X1 XNOR_1_1_NUM121 (.ZN (XNOR_1_1_NUM121_OUT), .A1 (N399), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM121 (.ZN (N447), .A1 (XNOR_1_1_NUM121_OUT), .A2 (GND));
      wire XNOR_1_1_NUM122_OUT;
      NOR2_X1 XNOR_1_1_NUM122 (.ZN (XNOR_1_1_NUM122_OUT), .A1 (N401), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM122 (.ZN (N448), .A1 (XNOR_1_1_NUM122_OUT), .A2 (GND));
      wire XNOR_1_1_NUM123_OUT;
      NOR2_X1 XNOR_1_1_NUM123 (.ZN (XNOR_1_1_NUM123_OUT), .A1 (N402), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM123 (.ZN (N449), .A1 (XNOR_1_1_NUM123_OUT), .A2 (GND));
      wire XNOR_1_1_NUM124_OUT;
      NOR2_X1 XNOR_1_1_NUM124 (.ZN (XNOR_1_1_NUM124_OUT), .A1 (N403), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM124 (.ZN (N450), .A1 (XNOR_1_1_NUM124_OUT), .A2 (GND));
      NOR2_X1 XNOR_NUM125 (.ZN (N451), .A1 (N424), .A2 (GND));
      NOR2_X1 XNOR_NUM126 (.ZN (N460), .A1 (N406), .A2 (N425));
      NOR2_X1 XNOR_NUM127 (.ZN (N463), .A1 (N409), .A2 (N426));
      wire XNOR_1_1_NUM128_OUT, XNOR_1_2_NUM128_OUT, XNOR_1_3_NUM128_OUT;
      NOR2_X1 XNOR_1_1_NUM128 (.ZN (XNOR_1_1_NUM128_OUT), .A1 (N442), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM128 (.ZN (XNOR_1_2_NUM128_OUT), .A1 (GND), .A2 (N410));
      NOR2_X1 XNOR_1_3_NUM128 (.ZN (XNOR_1_3_NUM128_OUT), .A1 (XNOR_1_1_NUM128_OUT), .A2 (XNOR_1_2_NUM128_OUT));
      NOR2_X1 XNOR_1_4_NUM128 (.ZN (N466), .A1 (XNOR_1_3_NUM128_OUT), .A2 (GND));
      wire XNOR_1_1_NUM129_OUT, XNOR_1_2_NUM129_OUT;
      NOR2_X1 XNOR_1_1_NUM129 (.ZN (XNOR_1_1_NUM129_OUT), .A1 (N143), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM129 (.ZN (XNOR_1_2_NUM129_OUT), .A1 (GND), .A2 (N427));
      NOR2_X1 XNOR_1_3_NUM129 (.ZN (N475), .A1 (XNOR_1_1_NUM129_OUT), .A2 (XNOR_1_2_NUM129_OUT));
      wire XNOR_1_1_NUM130_OUT, XNOR_1_2_NUM130_OUT;
      NOR2_X1 XNOR_1_1_NUM130 (.ZN (XNOR_1_1_NUM130_OUT), .A1 (N310), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM130 (.ZN (XNOR_1_2_NUM130_OUT), .A1 (GND), .A2 (N432));
      NOR2_X1 XNOR_1_3_NUM130 (.ZN (N476), .A1 (XNOR_1_1_NUM130_OUT), .A2 (XNOR_1_2_NUM130_OUT));
      wire XNOR_1_1_NUM131_OUT, XNOR_1_2_NUM131_OUT;
      NOR2_X1 XNOR_1_1_NUM131 (.ZN (XNOR_1_1_NUM131_OUT), .A1 (N146), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM131 (.ZN (XNOR_1_2_NUM131_OUT), .A1 (GND), .A2 (N427));
      NOR2_X1 XNOR_1_3_NUM131 (.ZN (N477), .A1 (XNOR_1_1_NUM131_OUT), .A2 (XNOR_1_2_NUM131_OUT));
      wire XNOR_1_1_NUM132_OUT, XNOR_1_2_NUM132_OUT;
      NOR2_X1 XNOR_1_1_NUM132 (.ZN (XNOR_1_1_NUM132_OUT), .A1 (N310), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM132 (.ZN (XNOR_1_2_NUM132_OUT), .A1 (GND), .A2 (N432));
      NOR2_X1 XNOR_1_3_NUM132 (.ZN (N478), .A1 (XNOR_1_1_NUM132_OUT), .A2 (XNOR_1_2_NUM132_OUT));
      wire XNOR_1_1_NUM133_OUT, XNOR_1_2_NUM133_OUT;
      NOR2_X1 XNOR_1_1_NUM133 (.ZN (XNOR_1_1_NUM133_OUT), .A1 (N149), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM133 (.ZN (XNOR_1_2_NUM133_OUT), .A1 (GND), .A2 (N427));
      NOR2_X1 XNOR_1_3_NUM133 (.ZN (N479), .A1 (XNOR_1_1_NUM133_OUT), .A2 (XNOR_1_2_NUM133_OUT));
      wire XNOR_1_1_NUM134_OUT, XNOR_1_2_NUM134_OUT;
      NOR2_X1 XNOR_1_1_NUM134 (.ZN (XNOR_1_1_NUM134_OUT), .A1 (N310), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM134 (.ZN (XNOR_1_2_NUM134_OUT), .A1 (GND), .A2 (N432));
      NOR2_X1 XNOR_1_3_NUM134 (.ZN (N480), .A1 (XNOR_1_1_NUM134_OUT), .A2 (XNOR_1_2_NUM134_OUT));
      wire XNOR_1_1_NUM135_OUT, XNOR_1_2_NUM135_OUT;
      NOR2_X1 XNOR_1_1_NUM135 (.ZN (XNOR_1_1_NUM135_OUT), .A1 (N153), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM135 (.ZN (XNOR_1_2_NUM135_OUT), .A1 (GND), .A2 (N427));
      NOR2_X1 XNOR_1_3_NUM135 (.ZN (N481), .A1 (XNOR_1_1_NUM135_OUT), .A2 (XNOR_1_2_NUM135_OUT));
      wire XNOR_1_1_NUM136_OUT, XNOR_1_2_NUM136_OUT;
      NOR2_X1 XNOR_1_1_NUM136 (.ZN (XNOR_1_1_NUM136_OUT), .A1 (N310), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM136 (.ZN (XNOR_1_2_NUM136_OUT), .A1 (GND), .A2 (N432));
      NOR2_X1 XNOR_1_3_NUM136 (.ZN (N482), .A1 (XNOR_1_1_NUM136_OUT), .A2 (XNOR_1_2_NUM136_OUT));
      wire XNOR_1_1_NUM137_OUT, XNOR_1_2_NUM137_OUT, XNOR_1_3_NUM137_OUT;
      NOR2_X1 XNOR_1_1_NUM137 (.ZN (XNOR_1_1_NUM137_OUT), .A1 (N443), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM137 (.ZN (XNOR_1_2_NUM137_OUT), .A1 (GND), .A2 (N1));
      NOR2_X1 XNOR_1_3_NUM137 (.ZN (XNOR_1_3_NUM137_OUT), .A1 (XNOR_1_1_NUM137_OUT), .A2 (XNOR_1_2_NUM137_OUT));
      NOR2_X1 XNOR_1_4_NUM137 (.ZN (N483), .A1 (XNOR_1_3_NUM137_OUT), .A2 (GND));
      wire XNOR_1_NUM138_OUT;
      NOR2_X1 XNOR_1_NUM138 (.ZN (XNOR_1_NUM138_OUT), .A1 (N369), .A2 (N437));
      NOR2_X1 XNOR_2_NUM138 (.ZN (N488), .A1 (XNOR_1_NUM138_OUT), .A2 (GND));
      wire XNOR_1_NUM139_OUT;
      NOR2_X1 XNOR_1_NUM139 (.ZN (XNOR_1_NUM139_OUT), .A1 (N369), .A2 (N437));
      NOR2_X1 XNOR_2_NUM139 (.ZN (N489), .A1 (XNOR_1_NUM139_OUT), .A2 (GND));
      wire XNOR_1_NUM140_OUT;
      NOR2_X1 XNOR_1_NUM140 (.ZN (XNOR_1_NUM140_OUT), .A1 (N369), .A2 (N437));
      NOR2_X1 XNOR_2_NUM140 (.ZN (N490), .A1 (XNOR_1_NUM140_OUT), .A2 (GND));
      wire XNOR_1_NUM141_OUT;
      NOR2_X1 XNOR_1_NUM141 (.ZN (XNOR_1_NUM141_OUT), .A1 (N369), .A2 (N437));
      NOR2_X1 XNOR_2_NUM141 (.ZN (N491), .A1 (XNOR_1_NUM141_OUT), .A2 (GND));
      NOR2_X1 XNOR_NUM142 (.ZN (N492), .A1 (N413), .A2 (N444));
      NOR2_X1 XNOR_NUM143 (.ZN (N495), .A1 (N416), .A2 (N445));
      wire XNOR_1_1_NUM144_OUT, XNOR_1_2_NUM144_OUT, XNOR_1_3_NUM144_OUT;
      NOR2_X1 XNOR_1_1_NUM144 (.ZN (XNOR_1_1_NUM144_OUT), .A1 (N130), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM144 (.ZN (XNOR_1_2_NUM144_OUT), .A1 (GND), .A2 (N460));
      NOR2_X1 XNOR_1_3_NUM144 (.ZN (XNOR_1_3_NUM144_OUT), .A1 (XNOR_1_1_NUM144_OUT), .A2 (XNOR_1_2_NUM144_OUT));
      NOR2_X1 XNOR_1_4_NUM144 (.ZN (N498), .A1 (XNOR_1_3_NUM144_OUT), .A2 (GND));
      wire XNOR_1_NUM145_OUT;
      NOR2_X1 XNOR_1_NUM145 (.ZN (XNOR_1_NUM145_OUT), .A1 (N130), .A2 (N460));
      NOR2_X1 XNOR_2_NUM145 (.ZN (N499), .A1 (XNOR_1_NUM145_OUT), .A2 (GND));
      wire XNOR_1_1_NUM146_OUT, XNOR_1_2_NUM146_OUT, XNOR_1_3_NUM146_OUT;
      NOR2_X1 XNOR_1_1_NUM146 (.ZN (XNOR_1_1_NUM146_OUT), .A1 (N463), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM146 (.ZN (XNOR_1_2_NUM146_OUT), .A1 (GND), .A2 (N135));
      NOR2_X1 XNOR_1_3_NUM146 (.ZN (XNOR_1_3_NUM146_OUT), .A1 (XNOR_1_1_NUM146_OUT), .A2 (XNOR_1_2_NUM146_OUT));
      NOR2_X1 XNOR_1_4_NUM146 (.ZN (N500), .A1 (XNOR_1_3_NUM146_OUT), .A2 (GND));
      wire XNOR_1_NUM147_OUT;
      NOR2_X1 XNOR_1_NUM147 (.ZN (XNOR_1_NUM147_OUT), .A1 (N463), .A2 (N135));
      NOR2_X1 XNOR_2_NUM147 (.ZN (N501), .A1 (XNOR_1_NUM147_OUT), .A2 (GND));
      wire XNOR_1_1_NUM148_OUT, XNOR_1_2_NUM148_OUT;
      NOR2_X1 XNOR_1_1_NUM148 (.ZN (XNOR_1_1_NUM148_OUT), .A1 (N91), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM148 (.ZN (XNOR_1_2_NUM148_OUT), .A1 (GND), .A2 (N466));
      NOR2_X1 XNOR_1_3_NUM148 (.ZN (N502), .A1 (XNOR_1_1_NUM148_OUT), .A2 (XNOR_1_2_NUM148_OUT));
      NOR2_X1 XNOR_NUM149 (.ZN (N503), .A1 (N475), .A2 (N476));
      wire XNOR_1_1_NUM150_OUT, XNOR_1_2_NUM150_OUT;
      NOR2_X1 XNOR_1_1_NUM150 (.ZN (XNOR_1_1_NUM150_OUT), .A1 (N96), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM150 (.ZN (XNOR_1_2_NUM150_OUT), .A1 (GND), .A2 (N466));
      NOR2_X1 XNOR_1_3_NUM150 (.ZN (N504), .A1 (XNOR_1_1_NUM150_OUT), .A2 (XNOR_1_2_NUM150_OUT));
      NOR2_X1 XNOR_NUM151 (.ZN (N505), .A1 (N477), .A2 (N478));
      wire XNOR_1_1_NUM152_OUT, XNOR_1_2_NUM152_OUT;
      NOR2_X1 XNOR_1_1_NUM152 (.ZN (XNOR_1_1_NUM152_OUT), .A1 (N101), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM152 (.ZN (XNOR_1_2_NUM152_OUT), .A1 (GND), .A2 (N466));
      NOR2_X1 XNOR_1_3_NUM152 (.ZN (N506), .A1 (XNOR_1_1_NUM152_OUT), .A2 (XNOR_1_2_NUM152_OUT));
      NOR2_X1 XNOR_NUM153 (.ZN (N507), .A1 (N479), .A2 (N480));
      wire XNOR_1_1_NUM154_OUT, XNOR_1_2_NUM154_OUT;
      NOR2_X1 XNOR_1_1_NUM154 (.ZN (XNOR_1_1_NUM154_OUT), .A1 (N106), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM154 (.ZN (XNOR_1_2_NUM154_OUT), .A1 (GND), .A2 (N466));
      NOR2_X1 XNOR_1_3_NUM154 (.ZN (N508), .A1 (XNOR_1_1_NUM154_OUT), .A2 (XNOR_1_2_NUM154_OUT));
      NOR2_X1 XNOR_NUM155 (.ZN (N509), .A1 (N481), .A2 (N482));
      wire XNOR_1_1_NUM156_OUT, XNOR_1_2_NUM156_OUT;
      NOR2_X1 XNOR_1_1_NUM156 (.ZN (XNOR_1_1_NUM156_OUT), .A1 (N143), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM156 (.ZN (XNOR_1_2_NUM156_OUT), .A1 (GND), .A2 (N483));
      NOR2_X1 XNOR_1_3_NUM156 (.ZN (N510), .A1 (XNOR_1_1_NUM156_OUT), .A2 (XNOR_1_2_NUM156_OUT));
      wire XNOR_1_1_NUM157_OUT, XNOR_1_2_NUM157_OUT;
      NOR2_X1 XNOR_1_1_NUM157 (.ZN (XNOR_1_1_NUM157_OUT), .A1 (N111), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM157 (.ZN (XNOR_1_2_NUM157_OUT), .A1 (GND), .A2 (N466));
      NOR2_X1 XNOR_1_3_NUM157 (.ZN (N511), .A1 (XNOR_1_1_NUM157_OUT), .A2 (XNOR_1_2_NUM157_OUT));
      wire XNOR_1_1_NUM158_OUT, XNOR_1_2_NUM158_OUT;
      NOR2_X1 XNOR_1_1_NUM158 (.ZN (XNOR_1_1_NUM158_OUT), .A1 (N146), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM158 (.ZN (XNOR_1_2_NUM158_OUT), .A1 (GND), .A2 (N483));
      NOR2_X1 XNOR_1_3_NUM158 (.ZN (N512), .A1 (XNOR_1_1_NUM158_OUT), .A2 (XNOR_1_2_NUM158_OUT));
      wire XNOR_1_1_NUM159_OUT, XNOR_1_2_NUM159_OUT;
      NOR2_X1 XNOR_1_1_NUM159 (.ZN (XNOR_1_1_NUM159_OUT), .A1 (N116), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM159 (.ZN (XNOR_1_2_NUM159_OUT), .A1 (GND), .A2 (N466));
      NOR2_X1 XNOR_1_3_NUM159 (.ZN (N513), .A1 (XNOR_1_1_NUM159_OUT), .A2 (XNOR_1_2_NUM159_OUT));
      wire XNOR_1_1_NUM160_OUT, XNOR_1_2_NUM160_OUT;
      NOR2_X1 XNOR_1_1_NUM160 (.ZN (XNOR_1_1_NUM160_OUT), .A1 (N149), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM160 (.ZN (XNOR_1_2_NUM160_OUT), .A1 (GND), .A2 (N483));
      NOR2_X1 XNOR_1_3_NUM160 (.ZN (N514), .A1 (XNOR_1_1_NUM160_OUT), .A2 (XNOR_1_2_NUM160_OUT));
      wire XNOR_1_1_NUM161_OUT, XNOR_1_2_NUM161_OUT;
      NOR2_X1 XNOR_1_1_NUM161 (.ZN (XNOR_1_1_NUM161_OUT), .A1 (N121), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM161 (.ZN (XNOR_1_2_NUM161_OUT), .A1 (GND), .A2 (N466));
      NOR2_X1 XNOR_1_3_NUM161 (.ZN (N515), .A1 (XNOR_1_1_NUM161_OUT), .A2 (XNOR_1_2_NUM161_OUT));
      wire XNOR_1_1_NUM162_OUT, XNOR_1_2_NUM162_OUT;
      NOR2_X1 XNOR_1_1_NUM162 (.ZN (XNOR_1_1_NUM162_OUT), .A1 (N153), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM162 (.ZN (XNOR_1_2_NUM162_OUT), .A1 (GND), .A2 (N483));
      NOR2_X1 XNOR_1_3_NUM162 (.ZN (N516), .A1 (XNOR_1_1_NUM162_OUT), .A2 (XNOR_1_2_NUM162_OUT));
      wire XNOR_1_1_NUM163_OUT, XNOR_1_2_NUM163_OUT;
      NOR2_X1 XNOR_1_1_NUM163 (.ZN (XNOR_1_1_NUM163_OUT), .A1 (N126), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM163 (.ZN (XNOR_1_2_NUM163_OUT), .A1 (GND), .A2 (N466));
      NOR2_X1 XNOR_1_3_NUM163 (.ZN (N517), .A1 (XNOR_1_1_NUM163_OUT), .A2 (XNOR_1_2_NUM163_OUT));
      wire XNOR_1_1_NUM164_OUT, XNOR_1_2_NUM164_OUT, XNOR_1_3_NUM164_OUT;
      NOR2_X1 XNOR_1_1_NUM164 (.ZN (XNOR_1_1_NUM164_OUT), .A1 (N130), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM164 (.ZN (XNOR_1_2_NUM164_OUT), .A1 (GND), .A2 (N492));
      NOR2_X1 XNOR_1_3_NUM164 (.ZN (XNOR_1_3_NUM164_OUT), .A1 (XNOR_1_1_NUM164_OUT), .A2 (XNOR_1_2_NUM164_OUT));
      NOR2_X1 XNOR_1_4_NUM164 (.ZN (N518), .A1 (XNOR_1_3_NUM164_OUT), .A2 (GND));
      wire XNOR_1_NUM165_OUT;
      NOR2_X1 XNOR_1_NUM165 (.ZN (XNOR_1_NUM165_OUT), .A1 (N130), .A2 (N492));
      NOR2_X1 XNOR_2_NUM165 (.ZN (N519), .A1 (XNOR_1_NUM165_OUT), .A2 (GND));
      wire XNOR_1_1_NUM166_OUT, XNOR_1_2_NUM166_OUT, XNOR_1_3_NUM166_OUT;
      NOR2_X1 XNOR_1_1_NUM166 (.ZN (XNOR_1_1_NUM166_OUT), .A1 (N495), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM166 (.ZN (XNOR_1_2_NUM166_OUT), .A1 (GND), .A2 (N207));
      NOR2_X1 XNOR_1_3_NUM166 (.ZN (XNOR_1_3_NUM166_OUT), .A1 (XNOR_1_1_NUM166_OUT), .A2 (XNOR_1_2_NUM166_OUT));
      NOR2_X1 XNOR_1_4_NUM166 (.ZN (N520), .A1 (XNOR_1_3_NUM166_OUT), .A2 (GND));
      wire XNOR_1_NUM167_OUT;
      NOR2_X1 XNOR_1_NUM167 (.ZN (XNOR_1_NUM167_OUT), .A1 (N495), .A2 (N207));
      NOR2_X1 XNOR_2_NUM167 (.ZN (N521), .A1 (XNOR_1_NUM167_OUT), .A2 (GND));
      wire XNOR_1_1_NUM168_OUT, XNOR_1_2_NUM168_OUT;
      NOR2_X1 XNOR_1_1_NUM168 (.ZN (XNOR_1_1_NUM168_OUT), .A1 (N451), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM168 (.ZN (XNOR_1_2_NUM168_OUT), .A1 (GND), .A2 (N159));
      NOR2_X1 XNOR_1_3_NUM168 (.ZN (N522), .A1 (XNOR_1_1_NUM168_OUT), .A2 (XNOR_1_2_NUM168_OUT));
      wire XNOR_1_1_NUM169_OUT, XNOR_1_2_NUM169_OUT;
      NOR2_X1 XNOR_1_1_NUM169 (.ZN (XNOR_1_1_NUM169_OUT), .A1 (N451), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM169 (.ZN (XNOR_1_2_NUM169_OUT), .A1 (GND), .A2 (N165));
      NOR2_X1 XNOR_1_3_NUM169 (.ZN (N523), .A1 (XNOR_1_1_NUM169_OUT), .A2 (XNOR_1_2_NUM169_OUT));
      wire XNOR_1_1_NUM170_OUT, XNOR_1_2_NUM170_OUT;
      NOR2_X1 XNOR_1_1_NUM170 (.ZN (XNOR_1_1_NUM170_OUT), .A1 (N451), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM170 (.ZN (XNOR_1_2_NUM170_OUT), .A1 (GND), .A2 (N171));
      NOR2_X1 XNOR_1_3_NUM170 (.ZN (N524), .A1 (XNOR_1_1_NUM170_OUT), .A2 (XNOR_1_2_NUM170_OUT));
      wire XNOR_1_1_NUM171_OUT, XNOR_1_2_NUM171_OUT;
      NOR2_X1 XNOR_1_1_NUM171 (.ZN (XNOR_1_1_NUM171_OUT), .A1 (N451), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM171 (.ZN (XNOR_1_2_NUM171_OUT), .A1 (GND), .A2 (N177));
      NOR2_X1 XNOR_1_3_NUM171 (.ZN (N525), .A1 (XNOR_1_1_NUM171_OUT), .A2 (XNOR_1_2_NUM171_OUT));
      wire XNOR_1_1_NUM172_OUT, XNOR_1_2_NUM172_OUT;
      NOR2_X1 XNOR_1_1_NUM172 (.ZN (XNOR_1_1_NUM172_OUT), .A1 (N451), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM172 (.ZN (XNOR_1_2_NUM172_OUT), .A1 (GND), .A2 (N183));
      NOR2_X1 XNOR_1_3_NUM172 (.ZN (N526), .A1 (XNOR_1_1_NUM172_OUT), .A2 (XNOR_1_2_NUM172_OUT));
      wire XNOR_1_1_NUM173_OUT, XNOR_1_2_NUM173_OUT, XNOR_1_3_NUM173_OUT;
      NOR2_X1 XNOR_1_1_NUM173 (.ZN (XNOR_1_1_NUM173_OUT), .A1 (N451), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM173 (.ZN (XNOR_1_2_NUM173_OUT), .A1 (GND), .A2 (N189));
      NOR2_X1 XNOR_1_3_NUM173 (.ZN (XNOR_1_3_NUM173_OUT), .A1 (XNOR_1_1_NUM173_OUT), .A2 (XNOR_1_2_NUM173_OUT));
      NOR2_X1 XNOR_1_4_NUM173 (.ZN (N527), .A1 (XNOR_1_3_NUM173_OUT), .A2 (GND));
      wire XNOR_1_1_NUM174_OUT, XNOR_1_2_NUM174_OUT, XNOR_1_3_NUM174_OUT;
      NOR2_X1 XNOR_1_1_NUM174 (.ZN (XNOR_1_1_NUM174_OUT), .A1 (N451), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM174 (.ZN (XNOR_1_2_NUM174_OUT), .A1 (GND), .A2 (N195));
      NOR2_X1 XNOR_1_3_NUM174 (.ZN (XNOR_1_3_NUM174_OUT), .A1 (XNOR_1_1_NUM174_OUT), .A2 (XNOR_1_2_NUM174_OUT));
      NOR2_X1 XNOR_1_4_NUM174 (.ZN (N528), .A1 (XNOR_1_3_NUM174_OUT), .A2 (GND));
      wire XNOR_1_1_NUM175_OUT, XNOR_1_2_NUM175_OUT, XNOR_1_3_NUM175_OUT;
      NOR2_X1 XNOR_1_1_NUM175 (.ZN (XNOR_1_1_NUM175_OUT), .A1 (N451), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM175 (.ZN (XNOR_1_2_NUM175_OUT), .A1 (GND), .A2 (N201));
      NOR2_X1 XNOR_1_3_NUM175 (.ZN (XNOR_1_3_NUM175_OUT), .A1 (XNOR_1_1_NUM175_OUT), .A2 (XNOR_1_2_NUM175_OUT));
      NOR2_X1 XNOR_1_4_NUM175 (.ZN (N529), .A1 (XNOR_1_3_NUM175_OUT), .A2 (GND));
      wire XNOR_1_1_NUM176_OUT, XNOR_1_2_NUM176_OUT, XNOR_1_3_NUM176_OUT;
      NOR2_X1 XNOR_1_1_NUM176 (.ZN (XNOR_1_1_NUM176_OUT), .A1 (N498), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM176 (.ZN (XNOR_1_2_NUM176_OUT), .A1 (GND), .A2 (N499));
      NOR2_X1 XNOR_1_3_NUM176 (.ZN (XNOR_1_3_NUM176_OUT), .A1 (XNOR_1_1_NUM176_OUT), .A2 (XNOR_1_2_NUM176_OUT));
      NOR2_X1 XNOR_1_4_NUM176 (.ZN (N530), .A1 (XNOR_1_3_NUM176_OUT), .A2 (GND));
      wire XNOR_1_1_NUM177_OUT, XNOR_1_2_NUM177_OUT, XNOR_1_3_NUM177_OUT;
      NOR2_X1 XNOR_1_1_NUM177 (.ZN (XNOR_1_1_NUM177_OUT), .A1 (N500), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM177 (.ZN (XNOR_1_2_NUM177_OUT), .A1 (GND), .A2 (N501));
      NOR2_X1 XNOR_1_3_NUM177 (.ZN (XNOR_1_3_NUM177_OUT), .A1 (XNOR_1_1_NUM177_OUT), .A2 (XNOR_1_2_NUM177_OUT));
      NOR2_X1 XNOR_1_4_NUM177 (.ZN (N533), .A1 (XNOR_1_3_NUM177_OUT), .A2 (GND));
      NOR2_X1 XNOR_NUM178 (.ZN (N536), .A1 (N309), .A2 (N502));
      NOR2_X1 XNOR_NUM179 (.ZN (N537), .A1 (N316), .A2 (N504));
      NOR2_X1 XNOR_NUM180 (.ZN (N538), .A1 (N317), .A2 (N506));
      NOR2_X1 XNOR_NUM181 (.ZN (N539), .A1 (N318), .A2 (N508));
      NOR2_X1 XNOR_NUM182 (.ZN (N540), .A1 (N510), .A2 (N511));
      NOR2_X1 XNOR_NUM183 (.ZN (N541), .A1 (N512), .A2 (N513));
      NOR2_X1 XNOR_NUM184 (.ZN (N542), .A1 (N514), .A2 (N515));
      NOR2_X1 XNOR_NUM185 (.ZN (N543), .A1 (N516), .A2 (N517));
      wire XNOR_1_1_NUM186_OUT, XNOR_1_2_NUM186_OUT, XNOR_1_3_NUM186_OUT;
      NOR2_X1 XNOR_1_1_NUM186 (.ZN (XNOR_1_1_NUM186_OUT), .A1 (N518), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM186 (.ZN (XNOR_1_2_NUM186_OUT), .A1 (GND), .A2 (N519));
      NOR2_X1 XNOR_1_3_NUM186 (.ZN (XNOR_1_3_NUM186_OUT), .A1 (XNOR_1_1_NUM186_OUT), .A2 (XNOR_1_2_NUM186_OUT));
      NOR2_X1 XNOR_1_4_NUM186 (.ZN (N544), .A1 (XNOR_1_3_NUM186_OUT), .A2 (GND));
      wire XNOR_1_1_NUM187_OUT, XNOR_1_2_NUM187_OUT, XNOR_1_3_NUM187_OUT;
      NOR2_X1 XNOR_1_1_NUM187 (.ZN (XNOR_1_1_NUM187_OUT), .A1 (N520), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM187 (.ZN (XNOR_1_2_NUM187_OUT), .A1 (GND), .A2 (N521));
      NOR2_X1 XNOR_1_3_NUM187 (.ZN (XNOR_1_3_NUM187_OUT), .A1 (XNOR_1_1_NUM187_OUT), .A2 (XNOR_1_2_NUM187_OUT));
      NOR2_X1 XNOR_1_4_NUM187 (.ZN (N547), .A1 (XNOR_1_3_NUM187_OUT), .A2 (GND));
      NOR2_X1 XNOR_NUM188 (.ZN (N550), .A1 (N530), .A2 (GND));
      NOR2_X1 XNOR_NUM189 (.ZN (N551), .A1 (N533), .A2 (GND));
      wire XNOR_1_1_NUM190_OUT, XNOR_1_2_NUM190_OUT;
      NOR2_X1 XNOR_1_1_NUM190 (.ZN (XNOR_1_1_NUM190_OUT), .A1 (N530), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM190 (.ZN (XNOR_1_2_NUM190_OUT), .A1 (GND), .A2 (N533));
      NOR2_X1 XNOR_1_3_NUM190 (.ZN (N552), .A1 (XNOR_1_1_NUM190_OUT), .A2 (XNOR_1_2_NUM190_OUT));
      wire XNOR_1_1_NUM191_OUT, XNOR_1_2_NUM191_OUT, XNOR_1_3_NUM191_OUT;
      NOR2_X1 XNOR_1_1_NUM191 (.ZN (XNOR_1_1_NUM191_OUT), .A1 (N536), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM191 (.ZN (XNOR_1_2_NUM191_OUT), .A1 (GND), .A2 (N503));
      NOR2_X1 XNOR_1_3_NUM191 (.ZN (XNOR_1_3_NUM191_OUT), .A1 (XNOR_1_1_NUM191_OUT), .A2 (XNOR_1_2_NUM191_OUT));
      NOR2_X1 XNOR_1_4_NUM191 (.ZN (N553), .A1 (XNOR_1_3_NUM191_OUT), .A2 (GND));
      wire XNOR_1_1_NUM192_OUT, XNOR_1_2_NUM192_OUT, XNOR_1_3_NUM192_OUT;
      NOR2_X1 XNOR_1_1_NUM192 (.ZN (XNOR_1_1_NUM192_OUT), .A1 (N537), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM192 (.ZN (XNOR_1_2_NUM192_OUT), .A1 (GND), .A2 (N505));
      NOR2_X1 XNOR_1_3_NUM192 (.ZN (XNOR_1_3_NUM192_OUT), .A1 (XNOR_1_1_NUM192_OUT), .A2 (XNOR_1_2_NUM192_OUT));
      NOR2_X1 XNOR_1_4_NUM192 (.ZN (N557), .A1 (XNOR_1_3_NUM192_OUT), .A2 (GND));
      wire XNOR_1_1_NUM193_OUT, XNOR_1_2_NUM193_OUT, XNOR_1_3_NUM193_OUT;
      NOR2_X1 XNOR_1_1_NUM193 (.ZN (XNOR_1_1_NUM193_OUT), .A1 (N538), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM193 (.ZN (XNOR_1_2_NUM193_OUT), .A1 (GND), .A2 (N507));
      NOR2_X1 XNOR_1_3_NUM193 (.ZN (XNOR_1_3_NUM193_OUT), .A1 (XNOR_1_1_NUM193_OUT), .A2 (XNOR_1_2_NUM193_OUT));
      NOR2_X1 XNOR_1_4_NUM193 (.ZN (N561), .A1 (XNOR_1_3_NUM193_OUT), .A2 (GND));
      wire XNOR_1_1_NUM194_OUT, XNOR_1_2_NUM194_OUT, XNOR_1_3_NUM194_OUT;
      NOR2_X1 XNOR_1_1_NUM194 (.ZN (XNOR_1_1_NUM194_OUT), .A1 (N539), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM194 (.ZN (XNOR_1_2_NUM194_OUT), .A1 (GND), .A2 (N509));
      NOR2_X1 XNOR_1_3_NUM194 (.ZN (XNOR_1_3_NUM194_OUT), .A1 (XNOR_1_1_NUM194_OUT), .A2 (XNOR_1_2_NUM194_OUT));
      NOR2_X1 XNOR_1_4_NUM194 (.ZN (N565), .A1 (XNOR_1_3_NUM194_OUT), .A2 (GND));
      wire XNOR_1_1_NUM195_OUT, XNOR_1_2_NUM195_OUT, XNOR_1_3_NUM195_OUT;
      NOR2_X1 XNOR_1_1_NUM195 (.ZN (XNOR_1_1_NUM195_OUT), .A1 (N488), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM195 (.ZN (XNOR_1_2_NUM195_OUT), .A1 (GND), .A2 (N540));
      NOR2_X1 XNOR_1_3_NUM195 (.ZN (XNOR_1_3_NUM195_OUT), .A1 (XNOR_1_1_NUM195_OUT), .A2 (XNOR_1_2_NUM195_OUT));
      NOR2_X1 XNOR_1_4_NUM195 (.ZN (N569), .A1 (XNOR_1_3_NUM195_OUT), .A2 (GND));
      wire XNOR_1_1_NUM196_OUT, XNOR_1_2_NUM196_OUT, XNOR_1_3_NUM196_OUT;
      NOR2_X1 XNOR_1_1_NUM196 (.ZN (XNOR_1_1_NUM196_OUT), .A1 (N489), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM196 (.ZN (XNOR_1_2_NUM196_OUT), .A1 (GND), .A2 (N541));
      NOR2_X1 XNOR_1_3_NUM196 (.ZN (XNOR_1_3_NUM196_OUT), .A1 (XNOR_1_1_NUM196_OUT), .A2 (XNOR_1_2_NUM196_OUT));
      NOR2_X1 XNOR_1_4_NUM196 (.ZN (N573), .A1 (XNOR_1_3_NUM196_OUT), .A2 (GND));
      wire XNOR_1_1_NUM197_OUT, XNOR_1_2_NUM197_OUT, XNOR_1_3_NUM197_OUT;
      NOR2_X1 XNOR_1_1_NUM197 (.ZN (XNOR_1_1_NUM197_OUT), .A1 (N490), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM197 (.ZN (XNOR_1_2_NUM197_OUT), .A1 (GND), .A2 (N542));
      NOR2_X1 XNOR_1_3_NUM197 (.ZN (XNOR_1_3_NUM197_OUT), .A1 (XNOR_1_1_NUM197_OUT), .A2 (XNOR_1_2_NUM197_OUT));
      NOR2_X1 XNOR_1_4_NUM197 (.ZN (N577), .A1 (XNOR_1_3_NUM197_OUT), .A2 (GND));
      wire XNOR_1_1_NUM198_OUT, XNOR_1_2_NUM198_OUT, XNOR_1_3_NUM198_OUT;
      NOR2_X1 XNOR_1_1_NUM198 (.ZN (XNOR_1_1_NUM198_OUT), .A1 (N491), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM198 (.ZN (XNOR_1_2_NUM198_OUT), .A1 (GND), .A2 (N543));
      NOR2_X1 XNOR_1_3_NUM198 (.ZN (XNOR_1_3_NUM198_OUT), .A1 (XNOR_1_1_NUM198_OUT), .A2 (XNOR_1_2_NUM198_OUT));
      NOR2_X1 XNOR_1_4_NUM198 (.ZN (N581), .A1 (XNOR_1_3_NUM198_OUT), .A2 (GND));
      NOR2_X1 XNOR_NUM199 (.ZN (N585), .A1 (N544), .A2 (GND));
      NOR2_X1 XNOR_NUM200 (.ZN (N586), .A1 (N547), .A2 (GND));
      wire XNOR_1_1_NUM201_OUT, XNOR_1_2_NUM201_OUT;
      NOR2_X1 XNOR_1_1_NUM201 (.ZN (XNOR_1_1_NUM201_OUT), .A1 (N544), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM201 (.ZN (XNOR_1_2_NUM201_OUT), .A1 (GND), .A2 (N547));
      NOR2_X1 XNOR_1_3_NUM201 (.ZN (N587), .A1 (XNOR_1_1_NUM201_OUT), .A2 (XNOR_1_2_NUM201_OUT));
      wire XNOR_1_1_NUM202_OUT, XNOR_1_2_NUM202_OUT;
      NOR2_X1 XNOR_1_1_NUM202 (.ZN (XNOR_1_1_NUM202_OUT), .A1 (N550), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM202 (.ZN (XNOR_1_2_NUM202_OUT), .A1 (GND), .A2 (N551));
      NOR2_X1 XNOR_1_3_NUM202 (.ZN (N588), .A1 (XNOR_1_1_NUM202_OUT), .A2 (XNOR_1_2_NUM202_OUT));
      wire XNOR_1_1_NUM203_OUT, XNOR_1_2_NUM203_OUT;
      NOR2_X1 XNOR_1_1_NUM203 (.ZN (XNOR_1_1_NUM203_OUT), .A1 (N585), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM203 (.ZN (XNOR_1_2_NUM203_OUT), .A1 (GND), .A2 (N586));
      NOR2_X1 XNOR_1_3_NUM203 (.ZN (N589), .A1 (XNOR_1_1_NUM203_OUT), .A2 (XNOR_1_2_NUM203_OUT));
      wire XNOR_1_1_NUM204_OUT, XNOR_1_2_NUM204_OUT, XNOR_1_3_NUM204_OUT;
      NOR2_X1 XNOR_1_1_NUM204 (.ZN (XNOR_1_1_NUM204_OUT), .A1 (N553), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM204 (.ZN (XNOR_1_2_NUM204_OUT), .A1 (GND), .A2 (N159));
      NOR2_X1 XNOR_1_3_NUM204 (.ZN (XNOR_1_3_NUM204_OUT), .A1 (XNOR_1_1_NUM204_OUT), .A2 (XNOR_1_2_NUM204_OUT));
      NOR2_X1 XNOR_1_4_NUM204 (.ZN (N590), .A1 (XNOR_1_3_NUM204_OUT), .A2 (GND));
      wire XNOR_1_NUM205_OUT;
      NOR2_X1 XNOR_1_NUM205 (.ZN (XNOR_1_NUM205_OUT), .A1 (N553), .A2 (N159));
      NOR2_X1 XNOR_2_NUM205 (.ZN (N593), .A1 (XNOR_1_NUM205_OUT), .A2 (GND));
      wire XNOR_1_1_NUM206_OUT, XNOR_1_2_NUM206_OUT;
      NOR2_X1 XNOR_1_1_NUM206 (.ZN (XNOR_1_1_NUM206_OUT), .A1 (N246), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM206 (.ZN (XNOR_1_2_NUM206_OUT), .A1 (GND), .A2 (N553));
      NOR2_X1 XNOR_1_3_NUM206 (.ZN (N596), .A1 (XNOR_1_1_NUM206_OUT), .A2 (XNOR_1_2_NUM206_OUT));
      wire XNOR_1_1_NUM207_OUT, XNOR_1_2_NUM207_OUT, XNOR_1_3_NUM207_OUT;
      NOR2_X1 XNOR_1_1_NUM207 (.ZN (XNOR_1_1_NUM207_OUT), .A1 (N557), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM207 (.ZN (XNOR_1_2_NUM207_OUT), .A1 (GND), .A2 (N165));
      NOR2_X1 XNOR_1_3_NUM207 (.ZN (XNOR_1_3_NUM207_OUT), .A1 (XNOR_1_1_NUM207_OUT), .A2 (XNOR_1_2_NUM207_OUT));
      NOR2_X1 XNOR_1_4_NUM207 (.ZN (N597), .A1 (XNOR_1_3_NUM207_OUT), .A2 (GND));
      wire XNOR_1_NUM208_OUT;
      NOR2_X1 XNOR_1_NUM208 (.ZN (XNOR_1_NUM208_OUT), .A1 (N557), .A2 (N165));
      NOR2_X1 XNOR_2_NUM208 (.ZN (N600), .A1 (XNOR_1_NUM208_OUT), .A2 (GND));
      wire XNOR_1_1_NUM209_OUT, XNOR_1_2_NUM209_OUT;
      NOR2_X1 XNOR_1_1_NUM209 (.ZN (XNOR_1_1_NUM209_OUT), .A1 (N246), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM209 (.ZN (XNOR_1_2_NUM209_OUT), .A1 (GND), .A2 (N557));
      NOR2_X1 XNOR_1_3_NUM209 (.ZN (N605), .A1 (XNOR_1_1_NUM209_OUT), .A2 (XNOR_1_2_NUM209_OUT));
      wire XNOR_1_1_NUM210_OUT, XNOR_1_2_NUM210_OUT, XNOR_1_3_NUM210_OUT;
      NOR2_X1 XNOR_1_1_NUM210 (.ZN (XNOR_1_1_NUM210_OUT), .A1 (N561), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM210 (.ZN (XNOR_1_2_NUM210_OUT), .A1 (GND), .A2 (N171));
      NOR2_X1 XNOR_1_3_NUM210 (.ZN (XNOR_1_3_NUM210_OUT), .A1 (XNOR_1_1_NUM210_OUT), .A2 (XNOR_1_2_NUM210_OUT));
      NOR2_X1 XNOR_1_4_NUM210 (.ZN (N606), .A1 (XNOR_1_3_NUM210_OUT), .A2 (GND));
      wire XNOR_1_NUM211_OUT;
      NOR2_X1 XNOR_1_NUM211 (.ZN (XNOR_1_NUM211_OUT), .A1 (N561), .A2 (N171));
      NOR2_X1 XNOR_2_NUM211 (.ZN (N609), .A1 (XNOR_1_NUM211_OUT), .A2 (GND));
      wire XNOR_1_1_NUM212_OUT, XNOR_1_2_NUM212_OUT;
      NOR2_X1 XNOR_1_1_NUM212 (.ZN (XNOR_1_1_NUM212_OUT), .A1 (N246), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM212 (.ZN (XNOR_1_2_NUM212_OUT), .A1 (GND), .A2 (N561));
      NOR2_X1 XNOR_1_3_NUM212 (.ZN (N615), .A1 (XNOR_1_1_NUM212_OUT), .A2 (XNOR_1_2_NUM212_OUT));
      wire XNOR_1_1_NUM213_OUT, XNOR_1_2_NUM213_OUT, XNOR_1_3_NUM213_OUT;
      NOR2_X1 XNOR_1_1_NUM213 (.ZN (XNOR_1_1_NUM213_OUT), .A1 (N565), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM213 (.ZN (XNOR_1_2_NUM213_OUT), .A1 (GND), .A2 (N177));
      NOR2_X1 XNOR_1_3_NUM213 (.ZN (XNOR_1_3_NUM213_OUT), .A1 (XNOR_1_1_NUM213_OUT), .A2 (XNOR_1_2_NUM213_OUT));
      NOR2_X1 XNOR_1_4_NUM213 (.ZN (N616), .A1 (XNOR_1_3_NUM213_OUT), .A2 (GND));
      wire XNOR_1_NUM214_OUT;
      NOR2_X1 XNOR_1_NUM214 (.ZN (XNOR_1_NUM214_OUT), .A1 (N565), .A2 (N177));
      NOR2_X1 XNOR_2_NUM214 (.ZN (N619), .A1 (XNOR_1_NUM214_OUT), .A2 (GND));
      wire XNOR_1_1_NUM215_OUT, XNOR_1_2_NUM215_OUT;
      NOR2_X1 XNOR_1_1_NUM215 (.ZN (XNOR_1_1_NUM215_OUT), .A1 (N246), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM215 (.ZN (XNOR_1_2_NUM215_OUT), .A1 (GND), .A2 (N565));
      NOR2_X1 XNOR_1_3_NUM215 (.ZN (N624), .A1 (XNOR_1_1_NUM215_OUT), .A2 (XNOR_1_2_NUM215_OUT));
      wire XNOR_1_1_NUM216_OUT, XNOR_1_2_NUM216_OUT, XNOR_1_3_NUM216_OUT;
      NOR2_X1 XNOR_1_1_NUM216 (.ZN (XNOR_1_1_NUM216_OUT), .A1 (N569), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM216 (.ZN (XNOR_1_2_NUM216_OUT), .A1 (GND), .A2 (N183));
      NOR2_X1 XNOR_1_3_NUM216 (.ZN (XNOR_1_3_NUM216_OUT), .A1 (XNOR_1_1_NUM216_OUT), .A2 (XNOR_1_2_NUM216_OUT));
      NOR2_X1 XNOR_1_4_NUM216 (.ZN (N625), .A1 (XNOR_1_3_NUM216_OUT), .A2 (GND));
      wire XNOR_1_NUM217_OUT;
      NOR2_X1 XNOR_1_NUM217 (.ZN (XNOR_1_NUM217_OUT), .A1 (N569), .A2 (N183));
      NOR2_X1 XNOR_2_NUM217 (.ZN (N628), .A1 (XNOR_1_NUM217_OUT), .A2 (GND));
      wire XNOR_1_1_NUM218_OUT, XNOR_1_2_NUM218_OUT;
      NOR2_X1 XNOR_1_1_NUM218 (.ZN (XNOR_1_1_NUM218_OUT), .A1 (N246), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM218 (.ZN (XNOR_1_2_NUM218_OUT), .A1 (GND), .A2 (N569));
      NOR2_X1 XNOR_1_3_NUM218 (.ZN (N631), .A1 (XNOR_1_1_NUM218_OUT), .A2 (XNOR_1_2_NUM218_OUT));
      wire XNOR_1_1_NUM219_OUT, XNOR_1_2_NUM219_OUT, XNOR_1_3_NUM219_OUT;
      NOR2_X1 XNOR_1_1_NUM219 (.ZN (XNOR_1_1_NUM219_OUT), .A1 (N573), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM219 (.ZN (XNOR_1_2_NUM219_OUT), .A1 (GND), .A2 (N189));
      NOR2_X1 XNOR_1_3_NUM219 (.ZN (XNOR_1_3_NUM219_OUT), .A1 (XNOR_1_1_NUM219_OUT), .A2 (XNOR_1_2_NUM219_OUT));
      NOR2_X1 XNOR_1_4_NUM219 (.ZN (N632), .A1 (XNOR_1_3_NUM219_OUT), .A2 (GND));
      wire XNOR_1_NUM220_OUT;
      NOR2_X1 XNOR_1_NUM220 (.ZN (XNOR_1_NUM220_OUT), .A1 (N573), .A2 (N189));
      NOR2_X1 XNOR_2_NUM220 (.ZN (N635), .A1 (XNOR_1_NUM220_OUT), .A2 (GND));
      wire XNOR_1_1_NUM221_OUT, XNOR_1_2_NUM221_OUT;
      NOR2_X1 XNOR_1_1_NUM221 (.ZN (XNOR_1_1_NUM221_OUT), .A1 (N246), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM221 (.ZN (XNOR_1_2_NUM221_OUT), .A1 (GND), .A2 (N573));
      NOR2_X1 XNOR_1_3_NUM221 (.ZN (N640), .A1 (XNOR_1_1_NUM221_OUT), .A2 (XNOR_1_2_NUM221_OUT));
      wire XNOR_1_1_NUM222_OUT, XNOR_1_2_NUM222_OUT, XNOR_1_3_NUM222_OUT;
      NOR2_X1 XNOR_1_1_NUM222 (.ZN (XNOR_1_1_NUM222_OUT), .A1 (N577), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM222 (.ZN (XNOR_1_2_NUM222_OUT), .A1 (GND), .A2 (N195));
      NOR2_X1 XNOR_1_3_NUM222 (.ZN (XNOR_1_3_NUM222_OUT), .A1 (XNOR_1_1_NUM222_OUT), .A2 (XNOR_1_2_NUM222_OUT));
      NOR2_X1 XNOR_1_4_NUM222 (.ZN (N641), .A1 (XNOR_1_3_NUM222_OUT), .A2 (GND));
      wire XNOR_1_NUM223_OUT;
      NOR2_X1 XNOR_1_NUM223 (.ZN (XNOR_1_NUM223_OUT), .A1 (N577), .A2 (N195));
      NOR2_X1 XNOR_2_NUM223 (.ZN (N644), .A1 (XNOR_1_NUM223_OUT), .A2 (GND));
      wire XNOR_1_1_NUM224_OUT, XNOR_1_2_NUM224_OUT;
      NOR2_X1 XNOR_1_1_NUM224 (.ZN (XNOR_1_1_NUM224_OUT), .A1 (N246), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM224 (.ZN (XNOR_1_2_NUM224_OUT), .A1 (GND), .A2 (N577));
      NOR2_X1 XNOR_1_3_NUM224 (.ZN (N650), .A1 (XNOR_1_1_NUM224_OUT), .A2 (XNOR_1_2_NUM224_OUT));
      wire XNOR_1_1_NUM225_OUT, XNOR_1_2_NUM225_OUT, XNOR_1_3_NUM225_OUT;
      NOR2_X1 XNOR_1_1_NUM225 (.ZN (XNOR_1_1_NUM225_OUT), .A1 (N581), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM225 (.ZN (XNOR_1_2_NUM225_OUT), .A1 (GND), .A2 (N201));
      NOR2_X1 XNOR_1_3_NUM225 (.ZN (XNOR_1_3_NUM225_OUT), .A1 (XNOR_1_1_NUM225_OUT), .A2 (XNOR_1_2_NUM225_OUT));
      NOR2_X1 XNOR_1_4_NUM225 (.ZN (N651), .A1 (XNOR_1_3_NUM225_OUT), .A2 (GND));
      wire XNOR_1_NUM226_OUT;
      NOR2_X1 XNOR_1_NUM226 (.ZN (XNOR_1_NUM226_OUT), .A1 (N581), .A2 (N201));
      NOR2_X1 XNOR_2_NUM226 (.ZN (N654), .A1 (XNOR_1_NUM226_OUT), .A2 (GND));
      wire XNOR_1_1_NUM227_OUT, XNOR_1_2_NUM227_OUT;
      NOR2_X1 XNOR_1_1_NUM227 (.ZN (XNOR_1_1_NUM227_OUT), .A1 (N246), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM227 (.ZN (XNOR_1_2_NUM227_OUT), .A1 (GND), .A2 (N581));
      NOR2_X1 XNOR_1_3_NUM227 (.ZN (N659), .A1 (XNOR_1_1_NUM227_OUT), .A2 (XNOR_1_2_NUM227_OUT));
      NOR2_X1 XNOR_NUM228 (.ZN (N660), .A1 (N552), .A2 (N588));
      NOR2_X1 XNOR_NUM229 (.ZN (N661), .A1 (N587), .A2 (N589));
      NOR2_X1 XNOR_NUM230 (.ZN (N662), .A1 (N590), .A2 (GND));
      wire XNOR_1_1_NUM231_OUT, XNOR_1_2_NUM231_OUT;
      NOR2_X1 XNOR_1_1_NUM231 (.ZN (XNOR_1_1_NUM231_OUT), .A1 (N593), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM231 (.ZN (XNOR_1_2_NUM231_OUT), .A1 (GND), .A2 (N590));
      NOR2_X1 XNOR_1_3_NUM231 (.ZN (N665), .A1 (XNOR_1_1_NUM231_OUT), .A2 (XNOR_1_2_NUM231_OUT));
      NOR2_X1 XNOR_NUM232 (.ZN (N669), .A1 (N596), .A2 (N522));
      NOR2_X1 XNOR_NUM233 (.ZN (N670), .A1 (N597), .A2 (GND));
      wire XNOR_1_1_NUM234_OUT, XNOR_1_2_NUM234_OUT;
      NOR2_X1 XNOR_1_1_NUM234 (.ZN (XNOR_1_1_NUM234_OUT), .A1 (N600), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM234 (.ZN (XNOR_1_2_NUM234_OUT), .A1 (GND), .A2 (N597));
      NOR2_X1 XNOR_1_3_NUM234 (.ZN (N673), .A1 (XNOR_1_1_NUM234_OUT), .A2 (XNOR_1_2_NUM234_OUT));
      NOR2_X1 XNOR_NUM235 (.ZN (N677), .A1 (N605), .A2 (N523));
      NOR2_X1 XNOR_NUM236 (.ZN (N678), .A1 (N606), .A2 (GND));
      wire XNOR_1_1_NUM237_OUT, XNOR_1_2_NUM237_OUT;
      NOR2_X1 XNOR_1_1_NUM237 (.ZN (XNOR_1_1_NUM237_OUT), .A1 (N609), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM237 (.ZN (XNOR_1_2_NUM237_OUT), .A1 (GND), .A2 (N606));
      NOR2_X1 XNOR_1_3_NUM237 (.ZN (N682), .A1 (XNOR_1_1_NUM237_OUT), .A2 (XNOR_1_2_NUM237_OUT));
      NOR2_X1 XNOR_NUM238 (.ZN (N686), .A1 (N615), .A2 (N524));
      NOR2_X1 XNOR_NUM239 (.ZN (N687), .A1 (N616), .A2 (GND));
      wire XNOR_1_1_NUM240_OUT, XNOR_1_2_NUM240_OUT;
      NOR2_X1 XNOR_1_1_NUM240 (.ZN (XNOR_1_1_NUM240_OUT), .A1 (N619), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM240 (.ZN (XNOR_1_2_NUM240_OUT), .A1 (GND), .A2 (N616));
      NOR2_X1 XNOR_1_3_NUM240 (.ZN (N692), .A1 (XNOR_1_1_NUM240_OUT), .A2 (XNOR_1_2_NUM240_OUT));
      NOR2_X1 XNOR_NUM241 (.ZN (N696), .A1 (N624), .A2 (N525));
      NOR2_X1 XNOR_NUM242 (.ZN (N697), .A1 (N625), .A2 (GND));
      wire XNOR_1_1_NUM243_OUT, XNOR_1_2_NUM243_OUT;
      NOR2_X1 XNOR_1_1_NUM243 (.ZN (XNOR_1_1_NUM243_OUT), .A1 (N628), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM243 (.ZN (XNOR_1_2_NUM243_OUT), .A1 (GND), .A2 (N625));
      NOR2_X1 XNOR_1_3_NUM243 (.ZN (N700), .A1 (XNOR_1_1_NUM243_OUT), .A2 (XNOR_1_2_NUM243_OUT));
      NOR2_X1 XNOR_NUM244 (.ZN (N704), .A1 (N631), .A2 (N526));
      NOR2_X1 XNOR_NUM245 (.ZN (N705), .A1 (N632), .A2 (GND));
      wire XNOR_1_1_NUM246_OUT, XNOR_1_2_NUM246_OUT;
      NOR2_X1 XNOR_1_1_NUM246 (.ZN (XNOR_1_1_NUM246_OUT), .A1 (N635), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM246 (.ZN (XNOR_1_2_NUM246_OUT), .A1 (GND), .A2 (N632));
      NOR2_X1 XNOR_1_3_NUM246 (.ZN (N708), .A1 (XNOR_1_1_NUM246_OUT), .A2 (XNOR_1_2_NUM246_OUT));
      NOR2_X1 XNOR_NUM247 (.ZN (N712), .A1 (N337), .A2 (N640));
      NOR2_X1 XNOR_NUM248 (.ZN (N713), .A1 (N641), .A2 (GND));
      wire XNOR_1_1_NUM249_OUT, XNOR_1_2_NUM249_OUT;
      NOR2_X1 XNOR_1_1_NUM249 (.ZN (XNOR_1_1_NUM249_OUT), .A1 (N644), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM249 (.ZN (XNOR_1_2_NUM249_OUT), .A1 (GND), .A2 (N641));
      NOR2_X1 XNOR_1_3_NUM249 (.ZN (N717), .A1 (XNOR_1_1_NUM249_OUT), .A2 (XNOR_1_2_NUM249_OUT));
      NOR2_X1 XNOR_NUM250 (.ZN (N721), .A1 (N339), .A2 (N650));
      NOR2_X1 XNOR_NUM251 (.ZN (N722), .A1 (N651), .A2 (GND));
      wire XNOR_1_1_NUM252_OUT, XNOR_1_2_NUM252_OUT;
      NOR2_X1 XNOR_1_1_NUM252 (.ZN (XNOR_1_1_NUM252_OUT), .A1 (N654), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM252 (.ZN (XNOR_1_2_NUM252_OUT), .A1 (GND), .A2 (N651));
      NOR2_X1 XNOR_1_3_NUM252 (.ZN (N727), .A1 (XNOR_1_1_NUM252_OUT), .A2 (XNOR_1_2_NUM252_OUT));
      NOR2_X1 XNOR_NUM253 (.ZN (N731), .A1 (N341), .A2 (N659));
      wire XNOR_1_1_NUM254_OUT, XNOR_1_2_NUM254_OUT, XNOR_1_3_NUM254_OUT;
      NOR2_X1 XNOR_1_1_NUM254 (.ZN (XNOR_1_1_NUM254_OUT), .A1 (N654), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM254 (.ZN (XNOR_1_2_NUM254_OUT), .A1 (GND), .A2 (N261));
      NOR2_X1 XNOR_1_3_NUM254 (.ZN (XNOR_1_3_NUM254_OUT), .A1 (XNOR_1_1_NUM254_OUT), .A2 (XNOR_1_2_NUM254_OUT));
      NOR2_X1 XNOR_1_4_NUM254 (.ZN (N732), .A1 (XNOR_1_3_NUM254_OUT), .A2 (GND));
      wire XNOR_1_1_NUM255_OUT, XNOR_1_2_NUM255_OUT, XNOR_1_3_NUM255_OUT;
      NOR2_X1 XNOR_1_1_NUM255 (.ZN (XNOR_1_1_NUM255_OUT), .A1 (N644), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM255 (.ZN (XNOR_1_2_NUM255_OUT), .A1 (GND), .A2 (N654));
      NOR2_X1 XNOR_1_3_NUM255 (.ZN (XNOR_1_3_NUM255_OUT), .A1 (XNOR_1_1_NUM255_OUT), .A2 (XNOR_1_2_NUM255_OUT));

      wire XNOR_2_1_NUM255_OUT, XNOR_2_2_NUM255_OUT, XNOR_2_3_NUM255_OUT;
      NOR2_X1 XNOR_2_1_NUM255 (.ZN (XNOR_2_1_NUM255_OUT), .A1 (N261), .A2 (GND));
      NOR2_X1 XNOR_2_2_NUM255 (.ZN (XNOR_2_2_NUM255_OUT), .A1 (GND), .A2 (XNOR_1_3_NUM255_OUT));
      NOR2_X1 XNOR_2_3_NUM255 (.ZN (XNOR_2_3_NUM255_OUT), .A1 (XNOR_2_1_NUM255_OUT), .A2 (XNOR_2_2_NUM255_OUT));

      NOR2_X1 XNOR_3_1_NUM255 (.ZN (N733), .A1 (XNOR_2_3_NUM255_OUT), .A2 (GND));
      wire XNOR_1_1_NUM256_OUT, XNOR_1_2_NUM256_OUT, XNOR_1_3_NUM256_OUT;
      NOR2_X1 XNOR_1_1_NUM256 (.ZN (XNOR_1_1_NUM256_OUT), .A1 (N635), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM256 (.ZN (XNOR_1_2_NUM256_OUT), .A1 (GND), .A2 (N644));
      NOR2_X1 XNOR_1_3_NUM256 (.ZN (XNOR_1_3_NUM256_OUT), .A1 (XNOR_1_1_NUM256_OUT), .A2 (XNOR_1_2_NUM256_OUT));

      wire XNOR_2_1_NUM256_OUT, XNOR_2_2_NUM256_OUT, XNOR_2_3_NUM256_OUT;
      NOR2_X1 XNOR_2_1_NUM256 (.ZN (XNOR_2_1_NUM256_OUT), .A1 (N654), .A2 (GND));
      NOR2_X1 XNOR_2_2_NUM256 (.ZN (XNOR_2_2_NUM256_OUT), .A1 (GND), .A2 (N261));
      NOR2_X1 XNOR_2_3_NUM256 (.ZN (XNOR_2_3_NUM256_OUT), .A1 (XNOR_2_1_NUM256_OUT), .A2 (XNOR_2_2_NUM256_OUT));

      wire XNOR_3_1_NUM256_OUT, XNOR_3_2_NUM256_OUT, XNOR_3_3_NUM256_OUT;
      NOR2_X1 XNOR_3_1_NUM256 (.ZN (XNOR_3_1_NUM256_OUT), .A1 (XNOR_1_3_NUM256_OUT), .A2 (GND));
      NOR2_X1 XNOR_3_2_NUM256 (.ZN (XNOR_3_2_NUM256_OUT), .A1 (GND), .A2 (XNOR_2_3_NUM256_OUT));
      NOR2_X1 XNOR_3_3_NUM256 (.ZN (XNOR_3_3_NUM256_OUT), .A1 (XNOR_3_1_NUM256_OUT), .A2 (XNOR_3_2_NUM256_OUT));

      NOR2_X1 XNOR_4_1_NUM256 (.ZN (N734), .A1 (XNOR_3_3_NUM256_OUT), .A2 (GND));
      NOR2_X1 XNOR_NUM257 (.ZN (N735), .A1 (N662), .A2 (GND));
      wire XNOR_1_1_NUM258_OUT, XNOR_1_2_NUM258_OUT;
      NOR2_X1 XNOR_1_1_NUM258 (.ZN (XNOR_1_1_NUM258_OUT), .A1 (N228), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM258 (.ZN (XNOR_1_2_NUM258_OUT), .A1 (GND), .A2 (N665));
      NOR2_X1 XNOR_1_3_NUM258 (.ZN (N736), .A1 (XNOR_1_1_NUM258_OUT), .A2 (XNOR_1_2_NUM258_OUT));
      wire XNOR_1_1_NUM259_OUT, XNOR_1_2_NUM259_OUT;
      NOR2_X1 XNOR_1_1_NUM259 (.ZN (XNOR_1_1_NUM259_OUT), .A1 (N237), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM259 (.ZN (XNOR_1_2_NUM259_OUT), .A1 (GND), .A2 (N662));
      NOR2_X1 XNOR_1_3_NUM259 (.ZN (N737), .A1 (XNOR_1_1_NUM259_OUT), .A2 (XNOR_1_2_NUM259_OUT));
      NOR2_X1 XNOR_NUM260 (.ZN (N738), .A1 (N670), .A2 (GND));
      wire XNOR_1_1_NUM261_OUT, XNOR_1_2_NUM261_OUT;
      NOR2_X1 XNOR_1_1_NUM261 (.ZN (XNOR_1_1_NUM261_OUT), .A1 (N228), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM261 (.ZN (XNOR_1_2_NUM261_OUT), .A1 (GND), .A2 (N673));
      NOR2_X1 XNOR_1_3_NUM261 (.ZN (N739), .A1 (XNOR_1_1_NUM261_OUT), .A2 (XNOR_1_2_NUM261_OUT));
      wire XNOR_1_1_NUM262_OUT, XNOR_1_2_NUM262_OUT;
      NOR2_X1 XNOR_1_1_NUM262 (.ZN (XNOR_1_1_NUM262_OUT), .A1 (N237), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM262 (.ZN (XNOR_1_2_NUM262_OUT), .A1 (GND), .A2 (N670));
      NOR2_X1 XNOR_1_3_NUM262 (.ZN (N740), .A1 (XNOR_1_1_NUM262_OUT), .A2 (XNOR_1_2_NUM262_OUT));
      NOR2_X1 XNOR_NUM263 (.ZN (N741), .A1 (N678), .A2 (GND));
      wire XNOR_1_1_NUM264_OUT, XNOR_1_2_NUM264_OUT;
      NOR2_X1 XNOR_1_1_NUM264 (.ZN (XNOR_1_1_NUM264_OUT), .A1 (N228), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM264 (.ZN (XNOR_1_2_NUM264_OUT), .A1 (GND), .A2 (N682));
      NOR2_X1 XNOR_1_3_NUM264 (.ZN (N742), .A1 (XNOR_1_1_NUM264_OUT), .A2 (XNOR_1_2_NUM264_OUT));
      wire XNOR_1_1_NUM265_OUT, XNOR_1_2_NUM265_OUT;
      NOR2_X1 XNOR_1_1_NUM265 (.ZN (XNOR_1_1_NUM265_OUT), .A1 (N237), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM265 (.ZN (XNOR_1_2_NUM265_OUT), .A1 (GND), .A2 (N678));
      NOR2_X1 XNOR_1_3_NUM265 (.ZN (N743), .A1 (XNOR_1_1_NUM265_OUT), .A2 (XNOR_1_2_NUM265_OUT));
      NOR2_X1 XNOR_NUM266 (.ZN (N744), .A1 (N687), .A2 (GND));
      wire XNOR_1_1_NUM267_OUT, XNOR_1_2_NUM267_OUT;
      NOR2_X1 XNOR_1_1_NUM267 (.ZN (XNOR_1_1_NUM267_OUT), .A1 (N228), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM267 (.ZN (XNOR_1_2_NUM267_OUT), .A1 (GND), .A2 (N692));
      NOR2_X1 XNOR_1_3_NUM267 (.ZN (N745), .A1 (XNOR_1_1_NUM267_OUT), .A2 (XNOR_1_2_NUM267_OUT));
      wire XNOR_1_1_NUM268_OUT, XNOR_1_2_NUM268_OUT;
      NOR2_X1 XNOR_1_1_NUM268 (.ZN (XNOR_1_1_NUM268_OUT), .A1 (N237), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM268 (.ZN (XNOR_1_2_NUM268_OUT), .A1 (GND), .A2 (N687));
      NOR2_X1 XNOR_1_3_NUM268 (.ZN (N746), .A1 (XNOR_1_1_NUM268_OUT), .A2 (XNOR_1_2_NUM268_OUT));
      NOR2_X1 XNOR_NUM269 (.ZN (N747), .A1 (N697), .A2 (GND));
      wire XNOR_1_1_NUM270_OUT, XNOR_1_2_NUM270_OUT;
      NOR2_X1 XNOR_1_1_NUM270 (.ZN (XNOR_1_1_NUM270_OUT), .A1 (N228), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM270 (.ZN (XNOR_1_2_NUM270_OUT), .A1 (GND), .A2 (N700));
      NOR2_X1 XNOR_1_3_NUM270 (.ZN (N748), .A1 (XNOR_1_1_NUM270_OUT), .A2 (XNOR_1_2_NUM270_OUT));
      wire XNOR_1_1_NUM271_OUT, XNOR_1_2_NUM271_OUT;
      NOR2_X1 XNOR_1_1_NUM271 (.ZN (XNOR_1_1_NUM271_OUT), .A1 (N237), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM271 (.ZN (XNOR_1_2_NUM271_OUT), .A1 (GND), .A2 (N697));
      NOR2_X1 XNOR_1_3_NUM271 (.ZN (N749), .A1 (XNOR_1_1_NUM271_OUT), .A2 (XNOR_1_2_NUM271_OUT));
      NOR2_X1 XNOR_NUM272 (.ZN (N750), .A1 (N705), .A2 (GND));
      wire XNOR_1_1_NUM273_OUT, XNOR_1_2_NUM273_OUT;
      NOR2_X1 XNOR_1_1_NUM273 (.ZN (XNOR_1_1_NUM273_OUT), .A1 (N228), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM273 (.ZN (XNOR_1_2_NUM273_OUT), .A1 (GND), .A2 (N708));
      NOR2_X1 XNOR_1_3_NUM273 (.ZN (N751), .A1 (XNOR_1_1_NUM273_OUT), .A2 (XNOR_1_2_NUM273_OUT));
      wire XNOR_1_1_NUM274_OUT, XNOR_1_2_NUM274_OUT;
      NOR2_X1 XNOR_1_1_NUM274 (.ZN (XNOR_1_1_NUM274_OUT), .A1 (N237), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM274 (.ZN (XNOR_1_2_NUM274_OUT), .A1 (GND), .A2 (N705));
      NOR2_X1 XNOR_1_3_NUM274 (.ZN (N752), .A1 (XNOR_1_1_NUM274_OUT), .A2 (XNOR_1_2_NUM274_OUT));
      NOR2_X1 XNOR_NUM275 (.ZN (N753), .A1 (N713), .A2 (GND));
      wire XNOR_1_1_NUM276_OUT, XNOR_1_2_NUM276_OUT;
      NOR2_X1 XNOR_1_1_NUM276 (.ZN (XNOR_1_1_NUM276_OUT), .A1 (N228), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM276 (.ZN (XNOR_1_2_NUM276_OUT), .A1 (GND), .A2 (N717));
      NOR2_X1 XNOR_1_3_NUM276 (.ZN (N754), .A1 (XNOR_1_1_NUM276_OUT), .A2 (XNOR_1_2_NUM276_OUT));
      wire XNOR_1_1_NUM277_OUT, XNOR_1_2_NUM277_OUT;
      NOR2_X1 XNOR_1_1_NUM277 (.ZN (XNOR_1_1_NUM277_OUT), .A1 (N237), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM277 (.ZN (XNOR_1_2_NUM277_OUT), .A1 (GND), .A2 (N713));
      NOR2_X1 XNOR_1_3_NUM277 (.ZN (N755), .A1 (XNOR_1_1_NUM277_OUT), .A2 (XNOR_1_2_NUM277_OUT));
      NOR2_X1 XNOR_NUM278 (.ZN (N756), .A1 (N722), .A2 (GND));
      NOR2_X1 XNOR_NUM279 (.ZN (N757), .A1 (N727), .A2 (N261));
      wire XNOR_1_1_NUM280_OUT, XNOR_1_2_NUM280_OUT;
      NOR2_X1 XNOR_1_1_NUM280 (.ZN (XNOR_1_1_NUM280_OUT), .A1 (N727), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM280 (.ZN (XNOR_1_2_NUM280_OUT), .A1 (GND), .A2 (N261));
      NOR2_X1 XNOR_1_3_NUM280 (.ZN (N758), .A1 (XNOR_1_1_NUM280_OUT), .A2 (XNOR_1_2_NUM280_OUT));
      wire XNOR_1_1_NUM281_OUT, XNOR_1_2_NUM281_OUT;
      NOR2_X1 XNOR_1_1_NUM281 (.ZN (XNOR_1_1_NUM281_OUT), .A1 (N228), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM281 (.ZN (XNOR_1_2_NUM281_OUT), .A1 (GND), .A2 (N727));
      NOR2_X1 XNOR_1_3_NUM281 (.ZN (N759), .A1 (XNOR_1_1_NUM281_OUT), .A2 (XNOR_1_2_NUM281_OUT));
      wire XNOR_1_1_NUM282_OUT, XNOR_1_2_NUM282_OUT;
      NOR2_X1 XNOR_1_1_NUM282 (.ZN (XNOR_1_1_NUM282_OUT), .A1 (N237), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM282 (.ZN (XNOR_1_2_NUM282_OUT), .A1 (GND), .A2 (N722));
      NOR2_X1 XNOR_1_3_NUM282 (.ZN (N760), .A1 (XNOR_1_1_NUM282_OUT), .A2 (XNOR_1_2_NUM282_OUT));
      wire XNOR_1_1_NUM283_OUT, XNOR_1_2_NUM283_OUT, XNOR_1_3_NUM283_OUT;
      NOR2_X1 XNOR_1_1_NUM283 (.ZN (XNOR_1_1_NUM283_OUT), .A1 (N644), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM283 (.ZN (XNOR_1_2_NUM283_OUT), .A1 (GND), .A2 (N722));
      NOR2_X1 XNOR_1_3_NUM283 (.ZN (XNOR_1_3_NUM283_OUT), .A1 (XNOR_1_1_NUM283_OUT), .A2 (XNOR_1_2_NUM283_OUT));
      NOR2_X1 XNOR_1_4_NUM283 (.ZN (N761), .A1 (XNOR_1_3_NUM283_OUT), .A2 (GND));
      wire XNOR_1_1_NUM284_OUT, XNOR_1_2_NUM284_OUT, XNOR_1_3_NUM284_OUT;
      NOR2_X1 XNOR_1_1_NUM284 (.ZN (XNOR_1_1_NUM284_OUT), .A1 (N635), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM284 (.ZN (XNOR_1_2_NUM284_OUT), .A1 (GND), .A2 (N713));
      NOR2_X1 XNOR_1_3_NUM284 (.ZN (XNOR_1_3_NUM284_OUT), .A1 (XNOR_1_1_NUM284_OUT), .A2 (XNOR_1_2_NUM284_OUT));
      NOR2_X1 XNOR_1_4_NUM284 (.ZN (N762), .A1 (XNOR_1_3_NUM284_OUT), .A2 (GND));
      wire XNOR_1_1_NUM285_OUT, XNOR_1_2_NUM285_OUT, XNOR_1_3_NUM285_OUT;
      NOR2_X1 XNOR_1_1_NUM285 (.ZN (XNOR_1_1_NUM285_OUT), .A1 (N635), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM285 (.ZN (XNOR_1_2_NUM285_OUT), .A1 (GND), .A2 (N644));
      NOR2_X1 XNOR_1_3_NUM285 (.ZN (XNOR_1_3_NUM285_OUT), .A1 (XNOR_1_1_NUM285_OUT), .A2 (XNOR_1_2_NUM285_OUT));

      wire XNOR_2_1_NUM285_OUT, XNOR_2_2_NUM285_OUT, XNOR_2_3_NUM285_OUT;
      NOR2_X1 XNOR_2_1_NUM285 (.ZN (XNOR_2_1_NUM285_OUT), .A1 (N722), .A2 (GND));
      NOR2_X1 XNOR_2_2_NUM285 (.ZN (XNOR_2_2_NUM285_OUT), .A1 (GND), .A2 (XNOR_1_3_NUM285_OUT));
      NOR2_X1 XNOR_2_3_NUM285 (.ZN (XNOR_2_3_NUM285_OUT), .A1 (XNOR_2_1_NUM285_OUT), .A2 (XNOR_2_2_NUM285_OUT));

      NOR2_X1 XNOR_3_1_NUM285 (.ZN (N763), .A1 (XNOR_2_3_NUM285_OUT), .A2 (GND));
      wire XNOR_1_1_NUM286_OUT, XNOR_1_2_NUM286_OUT, XNOR_1_3_NUM286_OUT;
      NOR2_X1 XNOR_1_1_NUM286 (.ZN (XNOR_1_1_NUM286_OUT), .A1 (N609), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM286 (.ZN (XNOR_1_2_NUM286_OUT), .A1 (GND), .A2 (N687));
      NOR2_X1 XNOR_1_3_NUM286 (.ZN (XNOR_1_3_NUM286_OUT), .A1 (XNOR_1_1_NUM286_OUT), .A2 (XNOR_1_2_NUM286_OUT));
      NOR2_X1 XNOR_1_4_NUM286 (.ZN (N764), .A1 (XNOR_1_3_NUM286_OUT), .A2 (GND));
      wire XNOR_1_1_NUM287_OUT, XNOR_1_2_NUM287_OUT, XNOR_1_3_NUM287_OUT;
      NOR2_X1 XNOR_1_1_NUM287 (.ZN (XNOR_1_1_NUM287_OUT), .A1 (N600), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM287 (.ZN (XNOR_1_2_NUM287_OUT), .A1 (GND), .A2 (N678));
      NOR2_X1 XNOR_1_3_NUM287 (.ZN (XNOR_1_3_NUM287_OUT), .A1 (XNOR_1_1_NUM287_OUT), .A2 (XNOR_1_2_NUM287_OUT));
      NOR2_X1 XNOR_1_4_NUM287 (.ZN (N765), .A1 (XNOR_1_3_NUM287_OUT), .A2 (GND));
      wire XNOR_1_1_NUM288_OUT, XNOR_1_2_NUM288_OUT, XNOR_1_3_NUM288_OUT;
      NOR2_X1 XNOR_1_1_NUM288 (.ZN (XNOR_1_1_NUM288_OUT), .A1 (N600), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM288 (.ZN (XNOR_1_2_NUM288_OUT), .A1 (GND), .A2 (N609));
      NOR2_X1 XNOR_1_3_NUM288 (.ZN (XNOR_1_3_NUM288_OUT), .A1 (XNOR_1_1_NUM288_OUT), .A2 (XNOR_1_2_NUM288_OUT));

      wire XNOR_2_1_NUM288_OUT, XNOR_2_2_NUM288_OUT, XNOR_2_3_NUM288_OUT;
      NOR2_X1 XNOR_2_1_NUM288 (.ZN (XNOR_2_1_NUM288_OUT), .A1 (N687), .A2 (GND));
      NOR2_X1 XNOR_2_2_NUM288 (.ZN (XNOR_2_2_NUM288_OUT), .A1 (GND), .A2 (XNOR_1_3_NUM288_OUT));
      NOR2_X1 XNOR_2_3_NUM288 (.ZN (XNOR_2_3_NUM288_OUT), .A1 (XNOR_2_1_NUM288_OUT), .A2 (XNOR_2_2_NUM288_OUT));

      NOR2_X1 XNOR_3_1_NUM288 (.ZN (N766), .A1 (XNOR_2_3_NUM288_OUT), .A2 (GND));
      wire XNOR_1_1_NUM289_OUT;
      NOR2_X1 XNOR_1_1_NUM289 (.ZN (XNOR_1_1_NUM289_OUT), .A1 (N660), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM289 (.ZN (N767), .A1 (XNOR_1_1_NUM289_OUT), .A2 (GND));
      wire XNOR_1_1_NUM290_OUT;
      NOR2_X1 XNOR_1_1_NUM290 (.ZN (XNOR_1_1_NUM290_OUT), .A1 (N661), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM290 (.ZN (N768), .A1 (XNOR_1_1_NUM290_OUT), .A2 (GND));
      NOR2_X1 XNOR_NUM291 (.ZN (N769), .A1 (N736), .A2 (N737));
      NOR2_X1 XNOR_NUM292 (.ZN (N770), .A1 (N739), .A2 (N740));
      NOR2_X1 XNOR_NUM293 (.ZN (N771), .A1 (N742), .A2 (N743));
      NOR2_X1 XNOR_NUM294 (.ZN (N772), .A1 (N745), .A2 (N746));
      wire XNOR_1_1_NUM295_OUT, XNOR_1_2_NUM295_OUT, XNOR_1_3_NUM295_OUT;
      NOR2_X1 XNOR_1_1_NUM295 (.ZN (XNOR_1_1_NUM295_OUT), .A1 (N750), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM295 (.ZN (XNOR_1_2_NUM295_OUT), .A1 (GND), .A2 (N762));
      NOR2_X1 XNOR_1_3_NUM295 (.ZN (XNOR_1_3_NUM295_OUT), .A1 (XNOR_1_1_NUM295_OUT), .A2 (XNOR_1_2_NUM295_OUT));

      wire XNOR_2_1_NUM295_OUT, XNOR_2_2_NUM295_OUT, XNOR_2_3_NUM295_OUT;
      NOR2_X1 XNOR_2_1_NUM295 (.ZN (XNOR_2_1_NUM295_OUT), .A1 (N763), .A2 (GND));
      NOR2_X1 XNOR_2_2_NUM295 (.ZN (XNOR_2_2_NUM295_OUT), .A1 (GND), .A2 (N734));
      NOR2_X1 XNOR_2_3_NUM295 (.ZN (XNOR_2_3_NUM295_OUT), .A1 (XNOR_2_1_NUM295_OUT), .A2 (XNOR_2_2_NUM295_OUT));

      wire XNOR_3_1_NUM295_OUT, XNOR_3_2_NUM295_OUT, XNOR_3_3_NUM295_OUT;
      NOR2_X1 XNOR_3_1_NUM295 (.ZN (XNOR_3_1_NUM295_OUT), .A1 (XNOR_1_3_NUM295_OUT), .A2 (GND));
      NOR2_X1 XNOR_3_2_NUM295 (.ZN (XNOR_3_2_NUM295_OUT), .A1 (GND), .A2 (XNOR_2_3_NUM295_OUT));
      NOR2_X1 XNOR_3_3_NUM295 (.ZN (XNOR_3_3_NUM295_OUT), .A1 (XNOR_3_1_NUM295_OUT), .A2 (XNOR_3_2_NUM295_OUT));

      NOR2_X1 XNOR_4_1_NUM295 (.ZN (N773), .A1 (XNOR_3_3_NUM295_OUT), .A2 (GND));
      NOR2_X1 XNOR_NUM296 (.ZN (N777), .A1 (N748), .A2 (N749));
      wire XNOR_1_1_NUM297_OUT, XNOR_1_2_NUM297_OUT, XNOR_1_3_NUM297_OUT;
      NOR2_X1 XNOR_1_1_NUM297 (.ZN (XNOR_1_1_NUM297_OUT), .A1 (N753), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM297 (.ZN (XNOR_1_2_NUM297_OUT), .A1 (GND), .A2 (N761));
      NOR2_X1 XNOR_1_3_NUM297 (.ZN (XNOR_1_3_NUM297_OUT), .A1 (XNOR_1_1_NUM297_OUT), .A2 (XNOR_1_2_NUM297_OUT));

      wire XNOR_2_1_NUM297_OUT, XNOR_2_2_NUM297_OUT, XNOR_2_3_NUM297_OUT;
      NOR2_X1 XNOR_2_1_NUM297 (.ZN (XNOR_2_1_NUM297_OUT), .A1 (N733), .A2 (GND));
      NOR2_X1 XNOR_2_2_NUM297 (.ZN (XNOR_2_2_NUM297_OUT), .A1 (GND), .A2 (XNOR_1_3_NUM297_OUT));
      NOR2_X1 XNOR_2_3_NUM297 (.ZN (XNOR_2_3_NUM297_OUT), .A1 (XNOR_2_1_NUM297_OUT), .A2 (XNOR_2_2_NUM297_OUT));

      NOR2_X1 XNOR_3_1_NUM297 (.ZN (N778), .A1 (XNOR_2_3_NUM297_OUT), .A2 (GND));
      NOR2_X1 XNOR_NUM298 (.ZN (N781), .A1 (N751), .A2 (N752));
      wire XNOR_1_1_NUM299_OUT, XNOR_1_2_NUM299_OUT, XNOR_1_3_NUM299_OUT;
      NOR2_X1 XNOR_1_1_NUM299 (.ZN (XNOR_1_1_NUM299_OUT), .A1 (N756), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM299 (.ZN (XNOR_1_2_NUM299_OUT), .A1 (GND), .A2 (N732));
      NOR2_X1 XNOR_1_3_NUM299 (.ZN (XNOR_1_3_NUM299_OUT), .A1 (XNOR_1_1_NUM299_OUT), .A2 (XNOR_1_2_NUM299_OUT));
      NOR2_X1 XNOR_1_4_NUM299 (.ZN (N782), .A1 (XNOR_1_3_NUM299_OUT), .A2 (GND));
      NOR2_X1 XNOR_NUM300 (.ZN (N785), .A1 (N754), .A2 (N755));
      NOR2_X1 XNOR_NUM301 (.ZN (N786), .A1 (N757), .A2 (N758));
      NOR2_X1 XNOR_NUM302 (.ZN (N787), .A1 (N759), .A2 (N760));
      NOR2_X1 XNOR_NUM303 (.ZN (N788), .A1 (N700), .A2 (N773));
      wire XNOR_1_1_NUM304_OUT, XNOR_1_2_NUM304_OUT;
      NOR2_X1 XNOR_1_1_NUM304 (.ZN (XNOR_1_1_NUM304_OUT), .A1 (N700), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM304 (.ZN (XNOR_1_2_NUM304_OUT), .A1 (GND), .A2 (N773));
      NOR2_X1 XNOR_1_3_NUM304 (.ZN (N789), .A1 (XNOR_1_1_NUM304_OUT), .A2 (XNOR_1_2_NUM304_OUT));
      NOR2_X1 XNOR_NUM305 (.ZN (N790), .A1 (N708), .A2 (N778));
      wire XNOR_1_1_NUM306_OUT, XNOR_1_2_NUM306_OUT;
      NOR2_X1 XNOR_1_1_NUM306 (.ZN (XNOR_1_1_NUM306_OUT), .A1 (N708), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM306 (.ZN (XNOR_1_2_NUM306_OUT), .A1 (GND), .A2 (N778));
      NOR2_X1 XNOR_1_3_NUM306 (.ZN (N791), .A1 (XNOR_1_1_NUM306_OUT), .A2 (XNOR_1_2_NUM306_OUT));
      NOR2_X1 XNOR_NUM307 (.ZN (N792), .A1 (N717), .A2 (N782));
      wire XNOR_1_1_NUM308_OUT, XNOR_1_2_NUM308_OUT;
      NOR2_X1 XNOR_1_1_NUM308 (.ZN (XNOR_1_1_NUM308_OUT), .A1 (N717), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM308 (.ZN (XNOR_1_2_NUM308_OUT), .A1 (GND), .A2 (N782));
      NOR2_X1 XNOR_1_3_NUM308 (.ZN (N793), .A1 (XNOR_1_1_NUM308_OUT), .A2 (XNOR_1_2_NUM308_OUT));
      wire XNOR_1_1_NUM309_OUT, XNOR_1_2_NUM309_OUT;
      NOR2_X1 XNOR_1_1_NUM309 (.ZN (XNOR_1_1_NUM309_OUT), .A1 (N219), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM309 (.ZN (XNOR_1_2_NUM309_OUT), .A1 (GND), .A2 (N786));
      NOR2_X1 XNOR_1_3_NUM309 (.ZN (N794), .A1 (XNOR_1_1_NUM309_OUT), .A2 (XNOR_1_2_NUM309_OUT));
      wire XNOR_1_1_NUM310_OUT, XNOR_1_2_NUM310_OUT, XNOR_1_3_NUM310_OUT;
      NOR2_X1 XNOR_1_1_NUM310 (.ZN (XNOR_1_1_NUM310_OUT), .A1 (N628), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM310 (.ZN (XNOR_1_2_NUM310_OUT), .A1 (GND), .A2 (N773));
      NOR2_X1 XNOR_1_3_NUM310 (.ZN (XNOR_1_3_NUM310_OUT), .A1 (XNOR_1_1_NUM310_OUT), .A2 (XNOR_1_2_NUM310_OUT));
      NOR2_X1 XNOR_1_4_NUM310 (.ZN (N795), .A1 (XNOR_1_3_NUM310_OUT), .A2 (GND));
      wire XNOR_1_1_NUM311_OUT, XNOR_1_2_NUM311_OUT, XNOR_1_3_NUM311_OUT;
      NOR2_X1 XNOR_1_1_NUM311 (.ZN (XNOR_1_1_NUM311_OUT), .A1 (N795), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM311 (.ZN (XNOR_1_2_NUM311_OUT), .A1 (GND), .A2 (N747));
      NOR2_X1 XNOR_1_3_NUM311 (.ZN (XNOR_1_3_NUM311_OUT), .A1 (XNOR_1_1_NUM311_OUT), .A2 (XNOR_1_2_NUM311_OUT));
      NOR2_X1 XNOR_1_4_NUM311 (.ZN (N796), .A1 (XNOR_1_3_NUM311_OUT), .A2 (GND));
      NOR2_X1 XNOR_NUM312 (.ZN (N802), .A1 (N788), .A2 (N789));
      NOR2_X1 XNOR_NUM313 (.ZN (N803), .A1 (N790), .A2 (N791));
      NOR2_X1 XNOR_NUM314 (.ZN (N804), .A1 (N792), .A2 (N793));
      NOR2_X1 XNOR_NUM315 (.ZN (N805), .A1 (N340), .A2 (N794));
      NOR2_X1 XNOR_NUM316 (.ZN (N806), .A1 (N692), .A2 (N796));
      wire XNOR_1_1_NUM317_OUT, XNOR_1_2_NUM317_OUT;
      NOR2_X1 XNOR_1_1_NUM317 (.ZN (XNOR_1_1_NUM317_OUT), .A1 (N692), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM317 (.ZN (XNOR_1_2_NUM317_OUT), .A1 (GND), .A2 (N796));
      NOR2_X1 XNOR_1_3_NUM317 (.ZN (N807), .A1 (XNOR_1_1_NUM317_OUT), .A2 (XNOR_1_2_NUM317_OUT));
      wire XNOR_1_1_NUM318_OUT, XNOR_1_2_NUM318_OUT;
      NOR2_X1 XNOR_1_1_NUM318 (.ZN (XNOR_1_1_NUM318_OUT), .A1 (N219), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM318 (.ZN (XNOR_1_2_NUM318_OUT), .A1 (GND), .A2 (N802));
      NOR2_X1 XNOR_1_3_NUM318 (.ZN (N808), .A1 (XNOR_1_1_NUM318_OUT), .A2 (XNOR_1_2_NUM318_OUT));
      wire XNOR_1_1_NUM319_OUT, XNOR_1_2_NUM319_OUT;
      NOR2_X1 XNOR_1_1_NUM319 (.ZN (XNOR_1_1_NUM319_OUT), .A1 (N219), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM319 (.ZN (XNOR_1_2_NUM319_OUT), .A1 (GND), .A2 (N803));
      NOR2_X1 XNOR_1_3_NUM319 (.ZN (N809), .A1 (XNOR_1_1_NUM319_OUT), .A2 (XNOR_1_2_NUM319_OUT));
      wire XNOR_1_1_NUM320_OUT, XNOR_1_2_NUM320_OUT;
      NOR2_X1 XNOR_1_1_NUM320 (.ZN (XNOR_1_1_NUM320_OUT), .A1 (N219), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM320 (.ZN (XNOR_1_2_NUM320_OUT), .A1 (GND), .A2 (N804));
      NOR2_X1 XNOR_1_3_NUM320 (.ZN (N810), .A1 (XNOR_1_1_NUM320_OUT), .A2 (XNOR_1_2_NUM320_OUT));
      wire XNOR_1_1_NUM321_OUT, XNOR_1_2_NUM321_OUT, XNOR_1_3_NUM321_OUT;
      NOR2_X1 XNOR_1_1_NUM321 (.ZN (XNOR_1_1_NUM321_OUT), .A1 (N805), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM321 (.ZN (XNOR_1_2_NUM321_OUT), .A1 (GND), .A2 (N787));
      NOR2_X1 XNOR_1_3_NUM321 (.ZN (XNOR_1_3_NUM321_OUT), .A1 (XNOR_1_1_NUM321_OUT), .A2 (XNOR_1_2_NUM321_OUT));

      wire XNOR_2_1_NUM321_OUT, XNOR_2_2_NUM321_OUT, XNOR_2_3_NUM321_OUT;
      NOR2_X1 XNOR_2_1_NUM321 (.ZN (XNOR_2_1_NUM321_OUT), .A1 (N731), .A2 (GND));
      NOR2_X1 XNOR_2_2_NUM321 (.ZN (XNOR_2_2_NUM321_OUT), .A1 (GND), .A2 (N529));
      NOR2_X1 XNOR_2_3_NUM321 (.ZN (XNOR_2_3_NUM321_OUT), .A1 (XNOR_2_1_NUM321_OUT), .A2 (XNOR_2_2_NUM321_OUT));

      wire XNOR_3_1_NUM321_OUT, XNOR_3_2_NUM321_OUT, XNOR_3_3_NUM321_OUT;
      NOR2_X1 XNOR_3_1_NUM321 (.ZN (XNOR_3_1_NUM321_OUT), .A1 (XNOR_1_3_NUM321_OUT), .A2 (GND));
      NOR2_X1 XNOR_3_2_NUM321 (.ZN (XNOR_3_2_NUM321_OUT), .A1 (GND), .A2 (XNOR_2_3_NUM321_OUT));
      NOR2_X1 XNOR_3_3_NUM321 (.ZN (XNOR_3_3_NUM321_OUT), .A1 (XNOR_3_1_NUM321_OUT), .A2 (XNOR_3_2_NUM321_OUT));

      NOR2_X1 XNOR_4_1_NUM321 (.ZN (N811), .A1 (XNOR_3_3_NUM321_OUT), .A2 (GND));
      wire XNOR_1_1_NUM322_OUT, XNOR_1_2_NUM322_OUT, XNOR_1_3_NUM322_OUT;
      NOR2_X1 XNOR_1_1_NUM322 (.ZN (XNOR_1_1_NUM322_OUT), .A1 (N619), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM322 (.ZN (XNOR_1_2_NUM322_OUT), .A1 (GND), .A2 (N796));
      NOR2_X1 XNOR_1_3_NUM322 (.ZN (XNOR_1_3_NUM322_OUT), .A1 (XNOR_1_1_NUM322_OUT), .A2 (XNOR_1_2_NUM322_OUT));
      NOR2_X1 XNOR_1_4_NUM322 (.ZN (N812), .A1 (XNOR_1_3_NUM322_OUT), .A2 (GND));
      wire XNOR_1_1_NUM323_OUT, XNOR_1_2_NUM323_OUT, XNOR_1_3_NUM323_OUT;
      NOR2_X1 XNOR_1_1_NUM323 (.ZN (XNOR_1_1_NUM323_OUT), .A1 (N609), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM323 (.ZN (XNOR_1_2_NUM323_OUT), .A1 (GND), .A2 (N619));
      NOR2_X1 XNOR_1_3_NUM323 (.ZN (XNOR_1_3_NUM323_OUT), .A1 (XNOR_1_1_NUM323_OUT), .A2 (XNOR_1_2_NUM323_OUT));

      wire XNOR_2_1_NUM323_OUT, XNOR_2_2_NUM323_OUT, XNOR_2_3_NUM323_OUT;
      NOR2_X1 XNOR_2_1_NUM323 (.ZN (XNOR_2_1_NUM323_OUT), .A1 (N796), .A2 (GND));
      NOR2_X1 XNOR_2_2_NUM323 (.ZN (XNOR_2_2_NUM323_OUT), .A1 (GND), .A2 (XNOR_1_3_NUM323_OUT));
      NOR2_X1 XNOR_2_3_NUM323 (.ZN (XNOR_2_3_NUM323_OUT), .A1 (XNOR_2_1_NUM323_OUT), .A2 (XNOR_2_2_NUM323_OUT));

      NOR2_X1 XNOR_3_1_NUM323 (.ZN (N813), .A1 (XNOR_2_3_NUM323_OUT), .A2 (GND));
      wire XNOR_1_1_NUM324_OUT, XNOR_1_2_NUM324_OUT, XNOR_1_3_NUM324_OUT;
      NOR2_X1 XNOR_1_1_NUM324 (.ZN (XNOR_1_1_NUM324_OUT), .A1 (N600), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM324 (.ZN (XNOR_1_2_NUM324_OUT), .A1 (GND), .A2 (N609));
      NOR2_X1 XNOR_1_3_NUM324 (.ZN (XNOR_1_3_NUM324_OUT), .A1 (XNOR_1_1_NUM324_OUT), .A2 (XNOR_1_2_NUM324_OUT));

      wire XNOR_2_1_NUM324_OUT, XNOR_2_2_NUM324_OUT, XNOR_2_3_NUM324_OUT;
      NOR2_X1 XNOR_2_1_NUM324 (.ZN (XNOR_2_1_NUM324_OUT), .A1 (N619), .A2 (GND));
      NOR2_X1 XNOR_2_2_NUM324 (.ZN (XNOR_2_2_NUM324_OUT), .A1 (GND), .A2 (N796));
      NOR2_X1 XNOR_2_3_NUM324 (.ZN (XNOR_2_3_NUM324_OUT), .A1 (XNOR_2_1_NUM324_OUT), .A2 (XNOR_2_2_NUM324_OUT));

      wire XNOR_3_1_NUM324_OUT, XNOR_3_2_NUM324_OUT, XNOR_3_3_NUM324_OUT;
      NOR2_X1 XNOR_3_1_NUM324 (.ZN (XNOR_3_1_NUM324_OUT), .A1 (XNOR_1_3_NUM324_OUT), .A2 (GND));
      NOR2_X1 XNOR_3_2_NUM324 (.ZN (XNOR_3_2_NUM324_OUT), .A1 (GND), .A2 (XNOR_2_3_NUM324_OUT));
      NOR2_X1 XNOR_3_3_NUM324 (.ZN (XNOR_3_3_NUM324_OUT), .A1 (XNOR_3_1_NUM324_OUT), .A2 (XNOR_3_2_NUM324_OUT));

      NOR2_X1 XNOR_4_1_NUM324 (.ZN (N814), .A1 (XNOR_3_3_NUM324_OUT), .A2 (GND));
      wire XNOR_1_1_NUM325_OUT, XNOR_1_2_NUM325_OUT, XNOR_1_3_NUM325_OUT;
      NOR2_X1 XNOR_1_1_NUM325 (.ZN (XNOR_1_1_NUM325_OUT), .A1 (N738), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM325 (.ZN (XNOR_1_2_NUM325_OUT), .A1 (GND), .A2 (N765));
      NOR2_X1 XNOR_1_3_NUM325 (.ZN (XNOR_1_3_NUM325_OUT), .A1 (XNOR_1_1_NUM325_OUT), .A2 (XNOR_1_2_NUM325_OUT));

      wire XNOR_2_1_NUM325_OUT, XNOR_2_2_NUM325_OUT, XNOR_2_3_NUM325_OUT;
      NOR2_X1 XNOR_2_1_NUM325 (.ZN (XNOR_2_1_NUM325_OUT), .A1 (N766), .A2 (GND));
      NOR2_X1 XNOR_2_2_NUM325 (.ZN (XNOR_2_2_NUM325_OUT), .A1 (GND), .A2 (N814));
      NOR2_X1 XNOR_2_3_NUM325 (.ZN (XNOR_2_3_NUM325_OUT), .A1 (XNOR_2_1_NUM325_OUT), .A2 (XNOR_2_2_NUM325_OUT));

      wire XNOR_3_1_NUM325_OUT, XNOR_3_2_NUM325_OUT, XNOR_3_3_NUM325_OUT;
      NOR2_X1 XNOR_3_1_NUM325 (.ZN (XNOR_3_1_NUM325_OUT), .A1 (XNOR_1_3_NUM325_OUT), .A2 (GND));
      NOR2_X1 XNOR_3_2_NUM325 (.ZN (XNOR_3_2_NUM325_OUT), .A1 (GND), .A2 (XNOR_2_3_NUM325_OUT));
      NOR2_X1 XNOR_3_3_NUM325 (.ZN (XNOR_3_3_NUM325_OUT), .A1 (XNOR_3_1_NUM325_OUT), .A2 (XNOR_3_2_NUM325_OUT));

      NOR2_X1 XNOR_4_1_NUM325 (.ZN (N815), .A1 (XNOR_3_3_NUM325_OUT), .A2 (GND));
      wire XNOR_1_1_NUM326_OUT, XNOR_1_2_NUM326_OUT, XNOR_1_3_NUM326_OUT;
      NOR2_X1 XNOR_1_1_NUM326 (.ZN (XNOR_1_1_NUM326_OUT), .A1 (N741), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM326 (.ZN (XNOR_1_2_NUM326_OUT), .A1 (GND), .A2 (N764));
      NOR2_X1 XNOR_1_3_NUM326 (.ZN (XNOR_1_3_NUM326_OUT), .A1 (XNOR_1_1_NUM326_OUT), .A2 (XNOR_1_2_NUM326_OUT));

      wire XNOR_2_1_NUM326_OUT, XNOR_2_2_NUM326_OUT, XNOR_2_3_NUM326_OUT;
      NOR2_X1 XNOR_2_1_NUM326 (.ZN (XNOR_2_1_NUM326_OUT), .A1 (N813), .A2 (GND));
      NOR2_X1 XNOR_2_2_NUM326 (.ZN (XNOR_2_2_NUM326_OUT), .A1 (GND), .A2 (XNOR_1_3_NUM326_OUT));
      NOR2_X1 XNOR_2_3_NUM326 (.ZN (XNOR_2_3_NUM326_OUT), .A1 (XNOR_2_1_NUM326_OUT), .A2 (XNOR_2_2_NUM326_OUT));

      NOR2_X1 XNOR_3_1_NUM326 (.ZN (N819), .A1 (XNOR_2_3_NUM326_OUT), .A2 (GND));
      wire XNOR_1_1_NUM327_OUT, XNOR_1_2_NUM327_OUT, XNOR_1_3_NUM327_OUT;
      NOR2_X1 XNOR_1_1_NUM327 (.ZN (XNOR_1_1_NUM327_OUT), .A1 (N744), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM327 (.ZN (XNOR_1_2_NUM327_OUT), .A1 (GND), .A2 (N812));
      NOR2_X1 XNOR_1_3_NUM327 (.ZN (XNOR_1_3_NUM327_OUT), .A1 (XNOR_1_1_NUM327_OUT), .A2 (XNOR_1_2_NUM327_OUT));
      NOR2_X1 XNOR_1_4_NUM327 (.ZN (N822), .A1 (XNOR_1_3_NUM327_OUT), .A2 (GND));
      NOR2_X1 XNOR_NUM328 (.ZN (N825), .A1 (N806), .A2 (N807));
      NOR2_X1 XNOR_NUM329 (.ZN (N826), .A1 (N335), .A2 (N808));
      NOR2_X1 XNOR_NUM330 (.ZN (N827), .A1 (N336), .A2 (N809));
      NOR2_X1 XNOR_NUM331 (.ZN (N828), .A1 (N338), .A2 (N810));
      NOR2_X1 XNOR_NUM332 (.ZN (N829), .A1 (N811), .A2 (GND));
      NOR2_X1 XNOR_NUM333 (.ZN (N830), .A1 (N665), .A2 (N815));
      wire XNOR_1_1_NUM334_OUT, XNOR_1_2_NUM334_OUT;
      NOR2_X1 XNOR_1_1_NUM334 (.ZN (XNOR_1_1_NUM334_OUT), .A1 (N665), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM334 (.ZN (XNOR_1_2_NUM334_OUT), .A1 (GND), .A2 (N815));
      NOR2_X1 XNOR_1_3_NUM334 (.ZN (N831), .A1 (XNOR_1_1_NUM334_OUT), .A2 (XNOR_1_2_NUM334_OUT));
      NOR2_X1 XNOR_NUM335 (.ZN (N832), .A1 (N673), .A2 (N819));
      wire XNOR_1_1_NUM336_OUT, XNOR_1_2_NUM336_OUT;
      NOR2_X1 XNOR_1_1_NUM336 (.ZN (XNOR_1_1_NUM336_OUT), .A1 (N673), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM336 (.ZN (XNOR_1_2_NUM336_OUT), .A1 (GND), .A2 (N819));
      NOR2_X1 XNOR_1_3_NUM336 (.ZN (N833), .A1 (XNOR_1_1_NUM336_OUT), .A2 (XNOR_1_2_NUM336_OUT));
      NOR2_X1 XNOR_NUM337 (.ZN (N834), .A1 (N682), .A2 (N822));
      wire XNOR_1_1_NUM338_OUT, XNOR_1_2_NUM338_OUT;
      NOR2_X1 XNOR_1_1_NUM338 (.ZN (XNOR_1_1_NUM338_OUT), .A1 (N682), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM338 (.ZN (XNOR_1_2_NUM338_OUT), .A1 (GND), .A2 (N822));
      NOR2_X1 XNOR_1_3_NUM338 (.ZN (N835), .A1 (XNOR_1_1_NUM338_OUT), .A2 (XNOR_1_2_NUM338_OUT));
      wire XNOR_1_1_NUM339_OUT, XNOR_1_2_NUM339_OUT;
      NOR2_X1 XNOR_1_1_NUM339 (.ZN (XNOR_1_1_NUM339_OUT), .A1 (N219), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM339 (.ZN (XNOR_1_2_NUM339_OUT), .A1 (GND), .A2 (N825));
      NOR2_X1 XNOR_1_3_NUM339 (.ZN (N836), .A1 (XNOR_1_1_NUM339_OUT), .A2 (XNOR_1_2_NUM339_OUT));
      wire XNOR_1_1_NUM340_OUT, XNOR_1_2_NUM340_OUT, XNOR_1_3_NUM340_OUT;
      NOR2_X1 XNOR_1_1_NUM340 (.ZN (XNOR_1_1_NUM340_OUT), .A1 (N826), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM340 (.ZN (XNOR_1_2_NUM340_OUT), .A1 (GND), .A2 (N777));
      NOR2_X1 XNOR_1_3_NUM340 (.ZN (XNOR_1_3_NUM340_OUT), .A1 (XNOR_1_1_NUM340_OUT), .A2 (XNOR_1_2_NUM340_OUT));

      wire XNOR_2_1_NUM340_OUT, XNOR_2_2_NUM340_OUT, XNOR_2_3_NUM340_OUT;
      NOR2_X1 XNOR_2_1_NUM340 (.ZN (XNOR_2_1_NUM340_OUT), .A1 (N704), .A2 (GND));
      NOR2_X1 XNOR_2_2_NUM340 (.ZN (XNOR_2_2_NUM340_OUT), .A1 (GND), .A2 (XNOR_1_3_NUM340_OUT));
      NOR2_X1 XNOR_2_3_NUM340 (.ZN (XNOR_2_3_NUM340_OUT), .A1 (XNOR_2_1_NUM340_OUT), .A2 (XNOR_2_2_NUM340_OUT));

      NOR2_X1 XNOR_3_1_NUM340 (.ZN (N837), .A1 (XNOR_2_3_NUM340_OUT), .A2 (GND));
      wire XNOR_1_1_NUM341_OUT, XNOR_1_2_NUM341_OUT, XNOR_1_3_NUM341_OUT;
      NOR2_X1 XNOR_1_1_NUM341 (.ZN (XNOR_1_1_NUM341_OUT), .A1 (N827), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM341 (.ZN (XNOR_1_2_NUM341_OUT), .A1 (GND), .A2 (N781));
      NOR2_X1 XNOR_1_3_NUM341 (.ZN (XNOR_1_3_NUM341_OUT), .A1 (XNOR_1_1_NUM341_OUT), .A2 (XNOR_1_2_NUM341_OUT));

      wire XNOR_2_1_NUM341_OUT, XNOR_2_2_NUM341_OUT, XNOR_2_3_NUM341_OUT;
      NOR2_X1 XNOR_2_1_NUM341 (.ZN (XNOR_2_1_NUM341_OUT), .A1 (N712), .A2 (GND));
      NOR2_X1 XNOR_2_2_NUM341 (.ZN (XNOR_2_2_NUM341_OUT), .A1 (GND), .A2 (N527));
      NOR2_X1 XNOR_2_3_NUM341 (.ZN (XNOR_2_3_NUM341_OUT), .A1 (XNOR_2_1_NUM341_OUT), .A2 (XNOR_2_2_NUM341_OUT));

      wire XNOR_3_1_NUM341_OUT, XNOR_3_2_NUM341_OUT, XNOR_3_3_NUM341_OUT;
      NOR2_X1 XNOR_3_1_NUM341 (.ZN (XNOR_3_1_NUM341_OUT), .A1 (XNOR_1_3_NUM341_OUT), .A2 (GND));
      NOR2_X1 XNOR_3_2_NUM341 (.ZN (XNOR_3_2_NUM341_OUT), .A1 (GND), .A2 (XNOR_2_3_NUM341_OUT));
      NOR2_X1 XNOR_3_3_NUM341 (.ZN (XNOR_3_3_NUM341_OUT), .A1 (XNOR_3_1_NUM341_OUT), .A2 (XNOR_3_2_NUM341_OUT));

      NOR2_X1 XNOR_4_1_NUM341 (.ZN (N838), .A1 (XNOR_3_3_NUM341_OUT), .A2 (GND));
      wire XNOR_1_1_NUM342_OUT, XNOR_1_2_NUM342_OUT, XNOR_1_3_NUM342_OUT;
      NOR2_X1 XNOR_1_1_NUM342 (.ZN (XNOR_1_1_NUM342_OUT), .A1 (N828), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM342 (.ZN (XNOR_1_2_NUM342_OUT), .A1 (GND), .A2 (N785));
      NOR2_X1 XNOR_1_3_NUM342 (.ZN (XNOR_1_3_NUM342_OUT), .A1 (XNOR_1_1_NUM342_OUT), .A2 (XNOR_1_2_NUM342_OUT));

      wire XNOR_2_1_NUM342_OUT, XNOR_2_2_NUM342_OUT, XNOR_2_3_NUM342_OUT;
      NOR2_X1 XNOR_2_1_NUM342 (.ZN (XNOR_2_1_NUM342_OUT), .A1 (N721), .A2 (GND));
      NOR2_X1 XNOR_2_2_NUM342 (.ZN (XNOR_2_2_NUM342_OUT), .A1 (GND), .A2 (N528));
      NOR2_X1 XNOR_2_3_NUM342 (.ZN (XNOR_2_3_NUM342_OUT), .A1 (XNOR_2_1_NUM342_OUT), .A2 (XNOR_2_2_NUM342_OUT));

      wire XNOR_3_1_NUM342_OUT, XNOR_3_2_NUM342_OUT, XNOR_3_3_NUM342_OUT;
      NOR2_X1 XNOR_3_1_NUM342 (.ZN (XNOR_3_1_NUM342_OUT), .A1 (XNOR_1_3_NUM342_OUT), .A2 (GND));
      NOR2_X1 XNOR_3_2_NUM342 (.ZN (XNOR_3_2_NUM342_OUT), .A1 (GND), .A2 (XNOR_2_3_NUM342_OUT));
      NOR2_X1 XNOR_3_3_NUM342 (.ZN (XNOR_3_3_NUM342_OUT), .A1 (XNOR_3_1_NUM342_OUT), .A2 (XNOR_3_2_NUM342_OUT));

      NOR2_X1 XNOR_4_1_NUM342 (.ZN (N839), .A1 (XNOR_3_3_NUM342_OUT), .A2 (GND));
      NOR2_X1 XNOR_NUM343 (.ZN (N840), .A1 (N829), .A2 (GND));
      wire XNOR_1_1_NUM344_OUT, XNOR_1_2_NUM344_OUT, XNOR_1_3_NUM344_OUT;
      NOR2_X1 XNOR_1_1_NUM344 (.ZN (XNOR_1_1_NUM344_OUT), .A1 (N815), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM344 (.ZN (XNOR_1_2_NUM344_OUT), .A1 (GND), .A2 (N593));
      NOR2_X1 XNOR_1_3_NUM344 (.ZN (XNOR_1_3_NUM344_OUT), .A1 (XNOR_1_1_NUM344_OUT), .A2 (XNOR_1_2_NUM344_OUT));
      NOR2_X1 XNOR_1_4_NUM344 (.ZN (N841), .A1 (XNOR_1_3_NUM344_OUT), .A2 (GND));
      NOR2_X1 XNOR_NUM345 (.ZN (N842), .A1 (N830), .A2 (N831));
      NOR2_X1 XNOR_NUM346 (.ZN (N843), .A1 (N832), .A2 (N833));
      NOR2_X1 XNOR_NUM347 (.ZN (N844), .A1 (N834), .A2 (N835));
      NOR2_X1 XNOR_NUM348 (.ZN (N845), .A1 (N334), .A2 (N836));
      NOR2_X1 XNOR_NUM349 (.ZN (N846), .A1 (N837), .A2 (GND));
      NOR2_X1 XNOR_NUM350 (.ZN (N847), .A1 (N838), .A2 (GND));
      NOR2_X1 XNOR_NUM351 (.ZN (N848), .A1 (N839), .A2 (GND));
      wire XNOR_1_1_NUM352_OUT, XNOR_1_2_NUM352_OUT;
      NOR2_X1 XNOR_1_1_NUM352 (.ZN (XNOR_1_1_NUM352_OUT), .A1 (N735), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM352 (.ZN (XNOR_1_2_NUM352_OUT), .A1 (GND), .A2 (N841));
      NOR2_X1 XNOR_1_3_NUM352 (.ZN (N849), .A1 (XNOR_1_1_NUM352_OUT), .A2 (XNOR_1_2_NUM352_OUT));
      wire XNOR_1_1_NUM353_OUT;
      NOR2_X1 XNOR_1_1_NUM353 (.ZN (XNOR_1_1_NUM353_OUT), .A1 (N840), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM353 (.ZN (N850), .A1 (XNOR_1_1_NUM353_OUT), .A2 (GND));
      wire XNOR_1_1_NUM354_OUT, XNOR_1_2_NUM354_OUT;
      NOR2_X1 XNOR_1_1_NUM354 (.ZN (XNOR_1_1_NUM354_OUT), .A1 (N219), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM354 (.ZN (XNOR_1_2_NUM354_OUT), .A1 (GND), .A2 (N842));
      NOR2_X1 XNOR_1_3_NUM354 (.ZN (N851), .A1 (XNOR_1_1_NUM354_OUT), .A2 (XNOR_1_2_NUM354_OUT));
      wire XNOR_1_1_NUM355_OUT, XNOR_1_2_NUM355_OUT;
      NOR2_X1 XNOR_1_1_NUM355 (.ZN (XNOR_1_1_NUM355_OUT), .A1 (N219), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM355 (.ZN (XNOR_1_2_NUM355_OUT), .A1 (GND), .A2 (N843));
      NOR2_X1 XNOR_1_3_NUM355 (.ZN (N852), .A1 (XNOR_1_1_NUM355_OUT), .A2 (XNOR_1_2_NUM355_OUT));
      wire XNOR_1_1_NUM356_OUT, XNOR_1_2_NUM356_OUT;
      NOR2_X1 XNOR_1_1_NUM356 (.ZN (XNOR_1_1_NUM356_OUT), .A1 (N219), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM356 (.ZN (XNOR_1_2_NUM356_OUT), .A1 (GND), .A2 (N844));
      NOR2_X1 XNOR_1_3_NUM356 (.ZN (N853), .A1 (XNOR_1_1_NUM356_OUT), .A2 (XNOR_1_2_NUM356_OUT));
      wire XNOR_1_1_NUM357_OUT, XNOR_1_2_NUM357_OUT, XNOR_1_3_NUM357_OUT;
      NOR2_X1 XNOR_1_1_NUM357 (.ZN (XNOR_1_1_NUM357_OUT), .A1 (N845), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM357 (.ZN (XNOR_1_2_NUM357_OUT), .A1 (GND), .A2 (N772));
      NOR2_X1 XNOR_1_3_NUM357 (.ZN (XNOR_1_3_NUM357_OUT), .A1 (XNOR_1_1_NUM357_OUT), .A2 (XNOR_1_2_NUM357_OUT));

      wire XNOR_2_1_NUM357_OUT, XNOR_2_2_NUM357_OUT, XNOR_2_3_NUM357_OUT;
      NOR2_X1 XNOR_2_1_NUM357 (.ZN (XNOR_2_1_NUM357_OUT), .A1 (N696), .A2 (GND));
      NOR2_X1 XNOR_2_2_NUM357 (.ZN (XNOR_2_2_NUM357_OUT), .A1 (GND), .A2 (XNOR_1_3_NUM357_OUT));
      NOR2_X1 XNOR_2_3_NUM357 (.ZN (XNOR_2_3_NUM357_OUT), .A1 (XNOR_2_1_NUM357_OUT), .A2 (XNOR_2_2_NUM357_OUT));

      NOR2_X1 XNOR_3_1_NUM357 (.ZN (N854), .A1 (XNOR_2_3_NUM357_OUT), .A2 (GND));
      NOR2_X1 XNOR_NUM358 (.ZN (N855), .A1 (N846), .A2 (GND));
      NOR2_X1 XNOR_NUM359 (.ZN (N856), .A1 (N847), .A2 (GND));
      NOR2_X1 XNOR_NUM360 (.ZN (N857), .A1 (N848), .A2 (GND));
      NOR2_X1 XNOR_NUM361 (.ZN (N858), .A1 (N849), .A2 (GND));
      NOR2_X1 XNOR_NUM362 (.ZN (N859), .A1 (N417), .A2 (N851));
      NOR2_X1 XNOR_NUM363 (.ZN (N860), .A1 (N332), .A2 (N852));
      NOR2_X1 XNOR_NUM364 (.ZN (N861), .A1 (N333), .A2 (N853));
      NOR2_X1 XNOR_NUM365 (.ZN (N862), .A1 (N854), .A2 (GND));
      wire XNOR_1_1_NUM366_OUT;
      NOR2_X1 XNOR_1_1_NUM366 (.ZN (XNOR_1_1_NUM366_OUT), .A1 (N855), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM366 (.ZN (N863), .A1 (XNOR_1_1_NUM366_OUT), .A2 (GND));
      wire XNOR_1_1_NUM367_OUT;
      NOR2_X1 XNOR_1_1_NUM367 (.ZN (XNOR_1_1_NUM367_OUT), .A1 (N856), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM367 (.ZN (N864), .A1 (XNOR_1_1_NUM367_OUT), .A2 (GND));
      wire XNOR_1_1_NUM368_OUT;
      NOR2_X1 XNOR_1_1_NUM368 (.ZN (XNOR_1_1_NUM368_OUT), .A1 (N857), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM368 (.ZN (N865), .A1 (XNOR_1_1_NUM368_OUT), .A2 (GND));
      wire XNOR_1_1_NUM369_OUT;
      NOR2_X1 XNOR_1_1_NUM369 (.ZN (XNOR_1_1_NUM369_OUT), .A1 (N858), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM369 (.ZN (N866), .A1 (XNOR_1_1_NUM369_OUT), .A2 (GND));
      wire XNOR_1_1_NUM370_OUT, XNOR_1_2_NUM370_OUT, XNOR_1_3_NUM370_OUT;
      NOR2_X1 XNOR_1_1_NUM370 (.ZN (XNOR_1_1_NUM370_OUT), .A1 (N859), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM370 (.ZN (XNOR_1_2_NUM370_OUT), .A1 (GND), .A2 (N769));
      NOR2_X1 XNOR_1_3_NUM370 (.ZN (XNOR_1_3_NUM370_OUT), .A1 (XNOR_1_1_NUM370_OUT), .A2 (XNOR_1_2_NUM370_OUT));

      wire XNOR_2_1_NUM370_OUT, XNOR_2_2_NUM370_OUT, XNOR_2_3_NUM370_OUT;
      NOR2_X1 XNOR_2_1_NUM370 (.ZN (XNOR_2_1_NUM370_OUT), .A1 (N669), .A2 (GND));
      NOR2_X1 XNOR_2_2_NUM370 (.ZN (XNOR_2_2_NUM370_OUT), .A1 (GND), .A2 (XNOR_1_3_NUM370_OUT));
      NOR2_X1 XNOR_2_3_NUM370 (.ZN (XNOR_2_3_NUM370_OUT), .A1 (XNOR_2_1_NUM370_OUT), .A2 (XNOR_2_2_NUM370_OUT));

      NOR2_X1 XNOR_3_1_NUM370 (.ZN (N867), .A1 (XNOR_2_3_NUM370_OUT), .A2 (GND));
      wire XNOR_1_1_NUM371_OUT, XNOR_1_2_NUM371_OUT, XNOR_1_3_NUM371_OUT;
      NOR2_X1 XNOR_1_1_NUM371 (.ZN (XNOR_1_1_NUM371_OUT), .A1 (N860), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM371 (.ZN (XNOR_1_2_NUM371_OUT), .A1 (GND), .A2 (N770));
      NOR2_X1 XNOR_1_3_NUM371 (.ZN (XNOR_1_3_NUM371_OUT), .A1 (XNOR_1_1_NUM371_OUT), .A2 (XNOR_1_2_NUM371_OUT));

      wire XNOR_2_1_NUM371_OUT, XNOR_2_2_NUM371_OUT, XNOR_2_3_NUM371_OUT;
      NOR2_X1 XNOR_2_1_NUM371 (.ZN (XNOR_2_1_NUM371_OUT), .A1 (N677), .A2 (GND));
      NOR2_X1 XNOR_2_2_NUM371 (.ZN (XNOR_2_2_NUM371_OUT), .A1 (GND), .A2 (XNOR_1_3_NUM371_OUT));
      NOR2_X1 XNOR_2_3_NUM371 (.ZN (XNOR_2_3_NUM371_OUT), .A1 (XNOR_2_1_NUM371_OUT), .A2 (XNOR_2_2_NUM371_OUT));

      NOR2_X1 XNOR_3_1_NUM371 (.ZN (N868), .A1 (XNOR_2_3_NUM371_OUT), .A2 (GND));
      wire XNOR_1_1_NUM372_OUT, XNOR_1_2_NUM372_OUT, XNOR_1_3_NUM372_OUT;
      NOR2_X1 XNOR_1_1_NUM372 (.ZN (XNOR_1_1_NUM372_OUT), .A1 (N861), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM372 (.ZN (XNOR_1_2_NUM372_OUT), .A1 (GND), .A2 (N771));
      NOR2_X1 XNOR_1_3_NUM372 (.ZN (XNOR_1_3_NUM372_OUT), .A1 (XNOR_1_1_NUM372_OUT), .A2 (XNOR_1_2_NUM372_OUT));

      wire XNOR_2_1_NUM372_OUT, XNOR_2_2_NUM372_OUT, XNOR_2_3_NUM372_OUT;
      NOR2_X1 XNOR_2_1_NUM372 (.ZN (XNOR_2_1_NUM372_OUT), .A1 (N686), .A2 (GND));
      NOR2_X1 XNOR_2_2_NUM372 (.ZN (XNOR_2_2_NUM372_OUT), .A1 (GND), .A2 (XNOR_1_3_NUM372_OUT));
      NOR2_X1 XNOR_2_3_NUM372 (.ZN (XNOR_2_3_NUM372_OUT), .A1 (XNOR_2_1_NUM372_OUT), .A2 (XNOR_2_2_NUM372_OUT));

      NOR2_X1 XNOR_3_1_NUM372 (.ZN (N869), .A1 (XNOR_2_3_NUM372_OUT), .A2 (GND));
      NOR2_X1 XNOR_NUM373 (.ZN (N870), .A1 (N862), .A2 (GND));
      NOR2_X1 XNOR_NUM374 (.ZN (N871), .A1 (N867), .A2 (GND));
      NOR2_X1 XNOR_NUM375 (.ZN (N872), .A1 (N868), .A2 (GND));
      NOR2_X1 XNOR_NUM376 (.ZN (N873), .A1 (N869), .A2 (GND));
      wire XNOR_1_1_NUM377_OUT;
      NOR2_X1 XNOR_1_1_NUM377 (.ZN (XNOR_1_1_NUM377_OUT), .A1 (N870), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM377 (.ZN (N874), .A1 (XNOR_1_1_NUM377_OUT), .A2 (GND));
      NOR2_X1 XNOR_NUM378 (.ZN (N875), .A1 (N871), .A2 (GND));
      NOR2_X1 XNOR_NUM379 (.ZN (N876), .A1 (N872), .A2 (GND));
      NOR2_X1 XNOR_NUM380 (.ZN (N877), .A1 (N873), .A2 (GND));
      wire XNOR_1_1_NUM381_OUT;
      NOR2_X1 XNOR_1_1_NUM381 (.ZN (XNOR_1_1_NUM381_OUT), .A1 (N875), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM381 (.ZN (N878), .A1 (XNOR_1_1_NUM381_OUT), .A2 (GND));
      wire XNOR_1_1_NUM382_OUT;
      NOR2_X1 XNOR_1_1_NUM382 (.ZN (XNOR_1_1_NUM382_OUT), .A1 (N876), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM382 (.ZN (N879), .A1 (XNOR_1_1_NUM382_OUT), .A2 (GND));
      wire XNOR_1_1_NUM383_OUT;
      NOR2_X1 XNOR_1_1_NUM383 (.ZN (XNOR_1_1_NUM383_OUT), .A1 (N877), .A2 (GND));
      NOR2_X1 XNOR_1_2_NUM383 (.ZN (N880), .A1 (XNOR_1_1_NUM383_OUT), .A2 (GND));


      wire XNOR_1_1_N388_TERMINATION_OUT, XNOR_1_2_N388_TERMINATION_OUT;
      NOR2_X1 XNOR_1_1_N388_TERMINATION (.ZN (XNOR_1_1_N388_TERMINATION_OUT), .A1 (N388), .A2 (GND));
      NOR2_X1 XNOR_1_2_N388_TERMINATION (.ZN (N388_TERMINATION), .A1 (XNOR_1_1_N388_TERMINATION_OUT), .A2 (XNOR_1_2_N388_TERMINATION_OUT));

      wire XNOR_1_1_N389_TERMINATION_OUT, XNOR_1_2_N389_TERMINATION_OUT;
      NOR2_X1 XNOR_1_1_N389_TERMINATION (.ZN (XNOR_1_1_N389_TERMINATION_OUT), .A1 (N389), .A2 (GND));
      NOR2_X1 XNOR_1_2_N389_TERMINATION (.ZN (N389_TERMINATION), .A1 (XNOR_1_1_N389_TERMINATION_OUT), .A2 (XNOR_1_2_N389_TERMINATION_OUT));

      wire XNOR_1_1_N390_TERMINATION_OUT, XNOR_1_2_N390_TERMINATION_OUT;
      NOR2_X1 XNOR_1_1_N390_TERMINATION (.ZN (XNOR_1_1_N390_TERMINATION_OUT), .A1 (N390), .A2 (GND));
      NOR2_X1 XNOR_1_2_N390_TERMINATION (.ZN (N390_TERMINATION), .A1 (XNOR_1_1_N390_TERMINATION_OUT), .A2 (XNOR_1_2_N390_TERMINATION_OUT));

      wire XNOR_1_1_N391_TERMINATION_OUT, XNOR_1_2_N391_TERMINATION_OUT;
      NOR2_X1 XNOR_1_1_N391_TERMINATION (.ZN (XNOR_1_1_N391_TERMINATION_OUT), .A1 (N391), .A2 (GND));
      NOR2_X1 XNOR_1_2_N391_TERMINATION (.ZN (N391_TERMINATION), .A1 (XNOR_1_1_N391_TERMINATION_OUT), .A2 (XNOR_1_2_N391_TERMINATION_OUT));

      wire XNOR_1_1_N418_TERMINATION_OUT, XNOR_1_2_N418_TERMINATION_OUT;
      NOR2_X1 XNOR_1_1_N418_TERMINATION (.ZN (XNOR_1_1_N418_TERMINATION_OUT), .A1 (N418), .A2 (GND));
      NOR2_X1 XNOR_1_2_N418_TERMINATION (.ZN (N418_TERMINATION), .A1 (XNOR_1_1_N418_TERMINATION_OUT), .A2 (XNOR_1_2_N418_TERMINATION_OUT));

      wire XNOR_1_1_N419_TERMINATION_OUT, XNOR_1_2_N419_TERMINATION_OUT;
      NOR2_X1 XNOR_1_1_N419_TERMINATION (.ZN (XNOR_1_1_N419_TERMINATION_OUT), .A1 (N419), .A2 (GND));
      NOR2_X1 XNOR_1_2_N419_TERMINATION (.ZN (N419_TERMINATION), .A1 (XNOR_1_1_N419_TERMINATION_OUT), .A2 (XNOR_1_2_N419_TERMINATION_OUT));

      wire XNOR_1_1_N420_TERMINATION_OUT, XNOR_1_2_N420_TERMINATION_OUT;
      NOR2_X1 XNOR_1_1_N420_TERMINATION (.ZN (XNOR_1_1_N420_TERMINATION_OUT), .A1 (N420), .A2 (GND));
      NOR2_X1 XNOR_1_2_N420_TERMINATION (.ZN (N420_TERMINATION), .A1 (XNOR_1_1_N420_TERMINATION_OUT), .A2 (XNOR_1_2_N420_TERMINATION_OUT));

      wire XNOR_1_1_N421_TERMINATION_OUT, XNOR_1_2_N421_TERMINATION_OUT;
      NOR2_X1 XNOR_1_1_N421_TERMINATION (.ZN (XNOR_1_1_N421_TERMINATION_OUT), .A1 (N421), .A2 (GND));
      NOR2_X1 XNOR_1_2_N421_TERMINATION (.ZN (N421_TERMINATION), .A1 (XNOR_1_1_N421_TERMINATION_OUT), .A2 (XNOR_1_2_N421_TERMINATION_OUT));

      wire XNOR_1_1_N422_TERMINATION_OUT, XNOR_1_2_N422_TERMINATION_OUT;
      NOR2_X1 XNOR_1_1_N422_TERMINATION (.ZN (XNOR_1_1_N422_TERMINATION_OUT), .A1 (N422), .A2 (GND));
      NOR2_X1 XNOR_1_2_N422_TERMINATION (.ZN (N422_TERMINATION), .A1 (XNOR_1_1_N422_TERMINATION_OUT), .A2 (XNOR_1_2_N422_TERMINATION_OUT));

      wire XNOR_1_1_N423_TERMINATION_OUT, XNOR_1_2_N423_TERMINATION_OUT;
      NOR2_X1 XNOR_1_1_N423_TERMINATION (.ZN (XNOR_1_1_N423_TERMINATION_OUT), .A1 (N423), .A2 (GND));
      NOR2_X1 XNOR_1_2_N423_TERMINATION (.ZN (N423_TERMINATION), .A1 (XNOR_1_1_N423_TERMINATION_OUT), .A2 (XNOR_1_2_N423_TERMINATION_OUT));

      wire XNOR_1_1_N446_TERMINATION_OUT, XNOR_1_2_N446_TERMINATION_OUT;
      NOR2_X1 XNOR_1_1_N446_TERMINATION (.ZN (XNOR_1_1_N446_TERMINATION_OUT), .A1 (N446), .A2 (GND));
      NOR2_X1 XNOR_1_2_N446_TERMINATION (.ZN (N446_TERMINATION), .A1 (XNOR_1_1_N446_TERMINATION_OUT), .A2 (XNOR_1_2_N446_TERMINATION_OUT));

      wire XNOR_1_1_N447_TERMINATION_OUT, XNOR_1_2_N447_TERMINATION_OUT;
      NOR2_X1 XNOR_1_1_N447_TERMINATION (.ZN (XNOR_1_1_N447_TERMINATION_OUT), .A1 (N447), .A2 (GND));
      NOR2_X1 XNOR_1_2_N447_TERMINATION (.ZN (N447_TERMINATION), .A1 (XNOR_1_1_N447_TERMINATION_OUT), .A2 (XNOR_1_2_N447_TERMINATION_OUT));

      wire XNOR_1_1_N448_TERMINATION_OUT, XNOR_1_2_N448_TERMINATION_OUT;
      NOR2_X1 XNOR_1_1_N448_TERMINATION (.ZN (XNOR_1_1_N448_TERMINATION_OUT), .A1 (N448), .A2 (GND));
      NOR2_X1 XNOR_1_2_N448_TERMINATION (.ZN (N448_TERMINATION), .A1 (XNOR_1_1_N448_TERMINATION_OUT), .A2 (XNOR_1_2_N448_TERMINATION_OUT));

      wire XNOR_1_1_N449_TERMINATION_OUT, XNOR_1_2_N449_TERMINATION_OUT;
      NOR2_X1 XNOR_1_1_N449_TERMINATION (.ZN (XNOR_1_1_N449_TERMINATION_OUT), .A1 (N449), .A2 (GND));
      NOR2_X1 XNOR_1_2_N449_TERMINATION (.ZN (N449_TERMINATION), .A1 (XNOR_1_1_N449_TERMINATION_OUT), .A2 (XNOR_1_2_N449_TERMINATION_OUT));

      wire XNOR_1_1_N450_TERMINATION_OUT, XNOR_1_2_N450_TERMINATION_OUT;
      NOR2_X1 XNOR_1_1_N450_TERMINATION (.ZN (XNOR_1_1_N450_TERMINATION_OUT), .A1 (N450), .A2 (GND));
      NOR2_X1 XNOR_1_2_N450_TERMINATION (.ZN (N450_TERMINATION), .A1 (XNOR_1_1_N450_TERMINATION_OUT), .A2 (XNOR_1_2_N450_TERMINATION_OUT));

      wire XNOR_1_1_N767_TERMINATION_OUT, XNOR_1_2_N767_TERMINATION_OUT;
      NOR2_X1 XNOR_1_1_N767_TERMINATION (.ZN (XNOR_1_1_N767_TERMINATION_OUT), .A1 (N767), .A2 (GND));
      NOR2_X1 XNOR_1_2_N767_TERMINATION (.ZN (N767_TERMINATION), .A1 (XNOR_1_1_N767_TERMINATION_OUT), .A2 (XNOR_1_2_N767_TERMINATION_OUT));

      wire XNOR_1_1_N768_TERMINATION_OUT, XNOR_1_2_N768_TERMINATION_OUT;
      NOR2_X1 XNOR_1_1_N768_TERMINATION (.ZN (XNOR_1_1_N768_TERMINATION_OUT), .A1 (N768), .A2 (GND));
      NOR2_X1 XNOR_1_2_N768_TERMINATION (.ZN (N768_TERMINATION), .A1 (XNOR_1_1_N768_TERMINATION_OUT), .A2 (XNOR_1_2_N768_TERMINATION_OUT));

      wire XNOR_1_1_N850_TERMINATION_OUT, XNOR_1_2_N850_TERMINATION_OUT;
      NOR2_X1 XNOR_1_1_N850_TERMINATION (.ZN (XNOR_1_1_N850_TERMINATION_OUT), .A1 (N850), .A2 (GND));
      NOR2_X1 XNOR_1_2_N850_TERMINATION (.ZN (N850_TERMINATION), .A1 (XNOR_1_1_N850_TERMINATION_OUT), .A2 (XNOR_1_2_N850_TERMINATION_OUT));

      wire XNOR_1_1_N863_TERMINATION_OUT, XNOR_1_2_N863_TERMINATION_OUT;
      NOR2_X1 XNOR_1_1_N863_TERMINATION (.ZN (XNOR_1_1_N863_TERMINATION_OUT), .A1 (N863), .A2 (GND));
      NOR2_X1 XNOR_1_2_N863_TERMINATION (.ZN (N863_TERMINATION), .A1 (XNOR_1_1_N863_TERMINATION_OUT), .A2 (XNOR_1_2_N863_TERMINATION_OUT));

      wire XNOR_1_1_N864_TERMINATION_OUT, XNOR_1_2_N864_TERMINATION_OUT;
      NOR2_X1 XNOR_1_1_N864_TERMINATION (.ZN (XNOR_1_1_N864_TERMINATION_OUT), .A1 (N864), .A2 (GND));
      NOR2_X1 XNOR_1_2_N864_TERMINATION (.ZN (N864_TERMINATION), .A1 (XNOR_1_1_N864_TERMINATION_OUT), .A2 (XNOR_1_2_N864_TERMINATION_OUT));

      wire XNOR_1_1_N865_TERMINATION_OUT, XNOR_1_2_N865_TERMINATION_OUT;
      NOR2_X1 XNOR_1_1_N865_TERMINATION (.ZN (XNOR_1_1_N865_TERMINATION_OUT), .A1 (N865), .A2 (GND));
      NOR2_X1 XNOR_1_2_N865_TERMINATION (.ZN (N865_TERMINATION), .A1 (XNOR_1_1_N865_TERMINATION_OUT), .A2 (XNOR_1_2_N865_TERMINATION_OUT));

      wire XNOR_1_1_N866_TERMINATION_OUT, XNOR_1_2_N866_TERMINATION_OUT;
      NOR2_X1 XNOR_1_1_N866_TERMINATION (.ZN (XNOR_1_1_N866_TERMINATION_OUT), .A1 (N866), .A2 (GND));
      NOR2_X1 XNOR_1_2_N866_TERMINATION (.ZN (N866_TERMINATION), .A1 (XNOR_1_1_N866_TERMINATION_OUT), .A2 (XNOR_1_2_N866_TERMINATION_OUT));

      wire XNOR_1_1_N874_TERMINATION_OUT, XNOR_1_2_N874_TERMINATION_OUT;
      NOR2_X1 XNOR_1_1_N874_TERMINATION (.ZN (XNOR_1_1_N874_TERMINATION_OUT), .A1 (N874), .A2 (GND));
      NOR2_X1 XNOR_1_2_N874_TERMINATION (.ZN (N874_TERMINATION), .A1 (XNOR_1_1_N874_TERMINATION_OUT), .A2 (XNOR_1_2_N874_TERMINATION_OUT));

      wire XNOR_1_1_N878_TERMINATION_OUT, XNOR_1_2_N878_TERMINATION_OUT;
      NOR2_X1 XNOR_1_1_N878_TERMINATION (.ZN (XNOR_1_1_N878_TERMINATION_OUT), .A1 (N878), .A2 (GND));
      NOR2_X1 XNOR_1_2_N878_TERMINATION (.ZN (N878_TERMINATION), .A1 (XNOR_1_1_N878_TERMINATION_OUT), .A2 (XNOR_1_2_N878_TERMINATION_OUT));

      wire XNOR_1_1_N879_TERMINATION_OUT, XNOR_1_2_N879_TERMINATION_OUT;
      NOR2_X1 XNOR_1_1_N879_TERMINATION (.ZN (XNOR_1_1_N879_TERMINATION_OUT), .A1 (N879), .A2 (GND));
      NOR2_X1 XNOR_1_2_N879_TERMINATION (.ZN (N879_TERMINATION), .A1 (XNOR_1_1_N879_TERMINATION_OUT), .A2 (XNOR_1_2_N879_TERMINATION_OUT));

      wire XNOR_1_1_N880_TERMINATION_OUT, XNOR_1_2_N880_TERMINATION_OUT;
      NOR2_X1 XNOR_1_1_N880_TERMINATION (.ZN (XNOR_1_1_N880_TERMINATION_OUT), .A1 (N880), .A2 (GND));
      NOR2_X1 XNOR_1_2_N880_TERMINATION (.ZN (N880_TERMINATION), .A1 (XNOR_1_1_N880_TERMINATION_OUT), .A2 (XNOR_1_2_N880_TERMINATION_OUT));


endmodule
* circuit: cgate_test
simulator lang=spice

*.PARAM pw=<sed>pw<sed>as
.PARAM supp=0.8V slope=0.1fs
.PARAM t_init0=0.1ns t_init1=0.174ns
.PARAM baseVal=0V peakVal=0.8V tend=2100.0ns


.LIB /home/s11777724/involution_tool_library_files/backend/spice/fet.inc CMG

* main circuit
.INCLUDE /home/s11777724/involution_tool_library_files/backend/spice/cell/BUF_X8.sp
.INCLUDE cgate.sp

**** SPECTRE Back Annotation
.option spef='/home/s11777724/JS/idm_evaluation/cgate_test/place_and_route/cgate_test_restitch.spef'
****

.TEMP 25
.OPTION
+ INGOLD=2
+ PARHIER=LOCAL
*+ POST=CSDF
+ PROBE
+ BRIEF
+ ACCURATE
+ ABSVAR=0.0001
+ DVDT=2
+ RELTOL=1e-11
*+ DELMAX=100fs
+ dc_pivot_check=yes

* vdd
VDD VDD GND 0.8v

.PARAM t_a_0=10ns
.PARAM t_a_1=13.333333ns
.PARAM t_a_2=15ns
.PARAM t_a_3=18.333333ns
.PARAM t_a_4=20ns
.PARAM t_a_5=23.333333ns
.PARAM t_a_6=25ns
.PARAM t_a_7=28.333333ns
.PARAM t_a_8=30ns
.PARAM t_a_9=33.333333ns
.PARAM t_a_10=35ns
.PARAM t_a_11=38.333333ns
.PARAM t_a_12=40ns
.PARAM t_a_13=43.333333ns
.PARAM t_a_14=45ns
.PARAM t_a_15=48.333333ns
.PARAM t_a_16=50ns
.PARAM t_a_17=53.333333ns
.PARAM t_a_18=55ns
.PARAM t_a_19=58.333333ns
.PARAM t_a_20=60ns
.PARAM t_a_21=63.333333ns
.PARAM t_a_22=65ns
.PARAM t_a_23=68.333333ns
.PARAM t_a_24=70ns
.PARAM t_a_25=73.333333ns
.PARAM t_a_26=75ns
.PARAM t_a_27=78.333333ns
.PARAM t_a_28=80ns
.PARAM t_a_29=83.333333ns
.PARAM t_a_30=85ns
.PARAM t_a_31=88.333333ns
.PARAM t_a_32=90ns
.PARAM t_a_33=93.333333ns
.PARAM t_a_34=95ns
.PARAM t_a_35=98.333333ns
.PARAM t_a_36=100ns
.PARAM t_a_37=103.333333ns
.PARAM t_a_38=105ns
.PARAM t_a_39=108.333333ns
.PARAM t_a_40=110ns
.PARAM t_a_41=113.333333ns
.PARAM t_a_42=115ns
.PARAM t_a_43=118.333333ns
.PARAM t_a_44=120ns
.PARAM t_a_45=123.333333ns
.PARAM t_a_46=125ns
.PARAM t_a_47=128.333333ns
.PARAM t_a_48=130ns
.PARAM t_a_49=133.333333ns
.PARAM t_a_50=135ns
.PARAM t_a_51=138.333333ns
.PARAM t_a_52=140ns
.PARAM t_a_53=143.333333ns
.PARAM t_a_54=145ns
.PARAM t_a_55=148.333333ns
.PARAM t_a_56=150ns
.PARAM t_a_57=153.333333ns
.PARAM t_a_58=155ns
.PARAM t_a_59=158.333333ns
.PARAM t_a_60=160ns
.PARAM t_a_61=163.333333ns
.PARAM t_a_62=165ns
.PARAM t_a_63=168.333333ns
.PARAM t_a_64=170ns
.PARAM t_a_65=173.333333ns
.PARAM t_a_66=175ns
.PARAM t_a_67=178.333333ns
.PARAM t_a_68=180ns
.PARAM t_a_69=183.333333ns
.PARAM t_a_70=185ns
.PARAM t_a_71=188.333333ns
.PARAM t_a_72=190ns
.PARAM t_a_73=193.333333ns
.PARAM t_a_74=195ns
.PARAM t_a_75=198.333333ns
.PARAM t_a_76=200ns
.PARAM t_a_77=203.333333ns
.PARAM t_a_78=205ns
.PARAM t_a_79=208.333333ns
.PARAM t_a_80=210ns
.PARAM t_a_81=213.333333ns
.PARAM t_a_82=215ns
.PARAM t_a_83=218.333333ns
.PARAM t_a_84=220ns
.PARAM t_a_85=223.333333ns
.PARAM t_a_86=225ns
.PARAM t_a_87=228.333333ns
.PARAM t_a_88=230ns
.PARAM t_a_89=233.333333ns
.PARAM t_a_90=235ns
.PARAM t_a_91=238.333333ns
.PARAM t_a_92=240ns
.PARAM t_a_93=243.333333ns
.PARAM t_a_94=245ns
.PARAM t_a_95=248.333333ns
.PARAM t_a_96=250ns
.PARAM t_a_97=253.333333ns
.PARAM t_a_98=255ns
.PARAM t_a_99=258.333333ns
.PARAM t_a_100=260ns
.PARAM t_a_101=263.333333ns
.PARAM t_a_102=265ns
.PARAM t_a_103=268.333333ns
.PARAM t_a_104=270ns
.PARAM t_a_105=273.333333ns
.PARAM t_a_106=275ns
.PARAM t_a_107=278.333333ns
.PARAM t_a_108=280ns
.PARAM t_a_109=283.333333ns
.PARAM t_a_110=285ns
.PARAM t_a_111=288.333333ns
.PARAM t_a_112=290ns
.PARAM t_a_113=293.333333ns
.PARAM t_a_114=295ns
.PARAM t_a_115=298.333333ns
.PARAM t_a_116=300ns
.PARAM t_a_117=303.333333ns
.PARAM t_a_118=305ns
.PARAM t_a_119=308.333333ns
.PARAM t_a_120=310ns
.PARAM t_a_121=313.333333ns
.PARAM t_a_122=315ns
.PARAM t_a_123=318.333333ns
.PARAM t_a_124=320ns
.PARAM t_a_125=323.333333ns
.PARAM t_a_126=325ns
.PARAM t_a_127=328.333333ns
.PARAM t_a_128=330ns
.PARAM t_a_129=333.333333ns
.PARAM t_a_130=335ns
.PARAM t_a_131=338.333333ns
.PARAM t_a_132=340ns
.PARAM t_a_133=343.333333ns
.PARAM t_a_134=345ns
.PARAM t_a_135=348.333333ns
.PARAM t_a_136=350ns
.PARAM t_a_137=353.333333ns
.PARAM t_a_138=355ns
.PARAM t_a_139=358.333333ns
.PARAM t_a_140=360ns
.PARAM t_a_141=363.333333ns
.PARAM t_a_142=365ns
.PARAM t_a_143=368.333333ns
.PARAM t_a_144=370ns
.PARAM t_a_145=373.333333ns
.PARAM t_a_146=375ns
.PARAM t_a_147=378.333333ns
.PARAM t_a_148=380ns
.PARAM t_a_149=383.333333ns
.PARAM t_a_150=385ns
.PARAM t_a_151=388.333333ns
.PARAM t_a_152=390ns
.PARAM t_a_153=393.333333ns
.PARAM t_a_154=395ns
.PARAM t_a_155=398.333333ns
.PARAM t_a_156=400ns
.PARAM t_a_157=403.333333ns
.PARAM t_a_158=405ns
.PARAM t_a_159=408.333333ns
.PARAM t_a_160=410ns
.PARAM t_a_161=413.333333ns
.PARAM t_a_162=415ns
.PARAM t_a_163=418.333333ns
.PARAM t_a_164=420ns
.PARAM t_a_165=423.333333ns
.PARAM t_a_166=425ns
.PARAM t_a_167=428.333333ns
.PARAM t_a_168=430ns
.PARAM t_a_169=433.333333ns
.PARAM t_a_170=435ns
.PARAM t_a_171=438.333333ns
.PARAM t_a_172=440ns
.PARAM t_a_173=443.333333ns
.PARAM t_a_174=445ns
.PARAM t_a_175=448.333333ns
.PARAM t_a_176=450ns
.PARAM t_a_177=453.333333ns
.PARAM t_a_178=455ns
.PARAM t_a_179=458.333333ns
.PARAM t_a_180=460ns
.PARAM t_a_181=463.333333ns
.PARAM t_a_182=465ns
.PARAM t_a_183=468.333333ns
.PARAM t_a_184=470ns
.PARAM t_a_185=473.333333ns
.PARAM t_a_186=475ns
.PARAM t_a_187=478.333333ns
.PARAM t_a_188=480ns
.PARAM t_a_189=483.333333ns
.PARAM t_a_190=485ns
.PARAM t_a_191=488.333333ns
.PARAM t_a_192=490ns
.PARAM t_a_193=493.333333ns
.PARAM t_a_194=495ns
.PARAM t_a_195=498.333333ns
.PARAM t_a_196=500ns
.PARAM t_a_197=503.333333ns
.PARAM t_a_198=505ns
.PARAM t_a_199=508.333333ns
.PARAM t_a_200=510ns
.PARAM t_a_201=513.333333ns
.PARAM t_a_202=515ns
.PARAM t_a_203=518.333333ns
.PARAM t_a_204=520ns
.PARAM t_a_205=523.333333ns
.PARAM t_a_206=525ns
.PARAM t_a_207=528.333333ns
.PARAM t_a_208=530ns
.PARAM t_a_209=533.333333ns
.PARAM t_a_210=535ns
.PARAM t_a_211=538.333333ns
.PARAM t_a_212=540ns
.PARAM t_a_213=543.333333ns
.PARAM t_a_214=545ns
.PARAM t_a_215=548.333333ns
.PARAM t_a_216=550ns
.PARAM t_a_217=553.333333ns
.PARAM t_a_218=555ns
.PARAM t_a_219=558.333333ns
.PARAM t_a_220=560ns
.PARAM t_a_221=563.333333ns
.PARAM t_a_222=565ns
.PARAM t_a_223=568.333333ns
.PARAM t_a_224=570ns
.PARAM t_a_225=573.333333ns
.PARAM t_a_226=575ns
.PARAM t_a_227=578.333333ns
.PARAM t_a_228=580ns
.PARAM t_a_229=583.333333ns
.PARAM t_a_230=585ns
.PARAM t_a_231=588.333333ns
.PARAM t_a_232=590ns
.PARAM t_a_233=593.333333ns
.PARAM t_a_234=595ns
.PARAM t_a_235=598.333333ns
.PARAM t_a_236=600ns
.PARAM t_a_237=603.333333ns
.PARAM t_a_238=605ns
.PARAM t_a_239=608.333333ns
.PARAM t_a_240=610ns
.PARAM t_a_241=613.333333ns
.PARAM t_a_242=615ns
.PARAM t_a_243=618.333333ns
.PARAM t_a_244=620ns
.PARAM t_a_245=623.333333ns
.PARAM t_a_246=625ns
.PARAM t_a_247=628.333333ns
.PARAM t_a_248=630ns
.PARAM t_a_249=633.333333ns
.PARAM t_a_250=635ns
.PARAM t_a_251=638.333333ns
.PARAM t_a_252=640ns
.PARAM t_a_253=643.333333ns
.PARAM t_a_254=645ns
.PARAM t_a_255=648.333333ns
.PARAM t_a_256=650ns
.PARAM t_a_257=653.333333ns
.PARAM t_a_258=655ns
.PARAM t_a_259=658.333333ns
.PARAM t_a_260=660ns
.PARAM t_a_261=663.333333ns
.PARAM t_a_262=665ns
.PARAM t_a_263=668.333333ns
.PARAM t_a_264=670ns
.PARAM t_a_265=673.333333ns
.PARAM t_a_266=675ns
.PARAM t_a_267=678.333333ns
.PARAM t_a_268=680ns
.PARAM t_a_269=683.333333ns
.PARAM t_a_270=685ns
.PARAM t_a_271=688.333333ns
.PARAM t_a_272=690ns
.PARAM t_a_273=693.333333ns
.PARAM t_a_274=695ns
.PARAM t_a_275=698.333333ns
.PARAM t_a_276=700ns
.PARAM t_a_277=703.333333ns
.PARAM t_a_278=705ns
.PARAM t_a_279=708.333333ns
.PARAM t_a_280=710ns
.PARAM t_a_281=713.333333ns
.PARAM t_a_282=715ns
.PARAM t_a_283=718.333333ns
.PARAM t_a_284=720ns
.PARAM t_a_285=723.333333ns
.PARAM t_a_286=725ns
.PARAM t_a_287=728.333333ns
.PARAM t_a_288=730ns
.PARAM t_a_289=733.333333ns
.PARAM t_a_290=735ns
.PARAM t_a_291=738.333333ns
.PARAM t_a_292=740ns
.PARAM t_a_293=743.333333ns
.PARAM t_a_294=745ns
.PARAM t_a_295=748.333333ns
.PARAM t_a_296=750ns
.PARAM t_a_297=753.333333ns
.PARAM t_a_298=755ns
.PARAM t_a_299=758.333333ns
.PARAM t_a_300=760ns
.PARAM t_a_301=763.333333ns
.PARAM t_a_302=765ns
.PARAM t_a_303=768.333333ns
.PARAM t_a_304=770ns
.PARAM t_a_305=773.333333ns
.PARAM t_a_306=775ns
.PARAM t_a_307=778.333333ns
.PARAM t_a_308=780ns
.PARAM t_a_309=783.333333ns
.PARAM t_a_310=785ns
.PARAM t_a_311=788.333333ns
.PARAM t_a_312=790ns
.PARAM t_a_313=793.333333ns
.PARAM t_a_314=795ns
.PARAM t_a_315=798.333333ns
.PARAM t_a_316=800ns
.PARAM t_a_317=803.333333ns
.PARAM t_a_318=805ns
.PARAM t_a_319=808.333333ns
.PARAM t_a_320=810ns
.PARAM t_a_321=813.333333ns
.PARAM t_a_322=815ns
.PARAM t_a_323=818.333333ns
.PARAM t_a_324=820ns
.PARAM t_a_325=823.333333ns
.PARAM t_a_326=825ns
.PARAM t_a_327=828.333333ns
.PARAM t_a_328=830ns
.PARAM t_a_329=833.333333ns
.PARAM t_a_330=835ns
.PARAM t_a_331=838.333333ns
.PARAM t_a_332=840ns
.PARAM t_a_333=843.333333ns
.PARAM t_a_334=845ns
.PARAM t_a_335=848.333333ns
.PARAM t_a_336=850ns
.PARAM t_a_337=853.333333ns
.PARAM t_a_338=855ns
.PARAM t_a_339=858.333333ns
.PARAM t_a_340=860ns
.PARAM t_a_341=863.333333ns
.PARAM t_a_342=865ns
.PARAM t_a_343=868.333333ns
.PARAM t_a_344=870ns
.PARAM t_a_345=873.333333ns
.PARAM t_a_346=875ns
.PARAM t_a_347=878.333333ns
.PARAM t_a_348=880ns
.PARAM t_a_349=883.333333ns
.PARAM t_a_350=885ns
.PARAM t_a_351=888.333333ns
.PARAM t_a_352=890ns
.PARAM t_a_353=893.333333ns
.PARAM t_a_354=895ns
.PARAM t_a_355=898.333333ns
.PARAM t_a_356=900ns
.PARAM t_a_357=903.333333ns
.PARAM t_a_358=905ns
.PARAM t_a_359=908.333333ns
.PARAM t_a_360=910ns
.PARAM t_a_361=913.333333ns
.PARAM t_a_362=915ns
.PARAM t_a_363=918.333333ns
.PARAM t_a_364=920ns
.PARAM t_a_365=923.333333ns
.PARAM t_a_366=925ns
.PARAM t_a_367=928.333333ns
.PARAM t_a_368=930ns
.PARAM t_a_369=933.333333ns
.PARAM t_a_370=935ns
.PARAM t_a_371=938.333333ns
.PARAM t_a_372=940ns
.PARAM t_a_373=943.333333ns
.PARAM t_a_374=945ns
.PARAM t_a_375=948.333333ns
.PARAM t_a_376=950ns
.PARAM t_a_377=953.333333ns
.PARAM t_a_378=955ns
.PARAM t_a_379=958.333333ns
.PARAM t_a_380=960ns
.PARAM t_a_381=963.333333ns
.PARAM t_a_382=965ns
.PARAM t_a_383=968.333333ns
.PARAM t_a_384=970ns
.PARAM t_a_385=973.333333ns
.PARAM t_a_386=975ns
.PARAM t_a_387=978.333333ns
.PARAM t_a_388=980ns
.PARAM t_a_389=983.333333ns
.PARAM t_a_390=985ns
.PARAM t_a_391=988.333333ns
.PARAM t_a_392=990ns
.PARAM t_a_393=993.333333ns
.PARAM t_a_394=995ns
.PARAM t_a_395=998.333333ns
.PARAM t_a_396=1000ns
.PARAM t_a_397=1003.333333ns
.PARAM t_a_398=1005ns
.PARAM t_a_399=1008.333333ns
.PARAM t_a_400=1010ns
.PARAM t_a_401=1013.333333ns
.PARAM t_a_402=1015ns
.PARAM t_a_403=1018.333333ns
.PARAM t_a_404=1020ns
.PARAM t_a_405=1023.333333ns
.PARAM t_a_406=1025ns
.PARAM t_a_407=1028.333333ns
.PARAM t_a_408=1030ns
.PARAM t_a_409=1033.333333ns
.PARAM t_a_410=1035ns
.PARAM t_a_411=1038.333333ns
.PARAM t_a_412=1040ns
.PARAM t_a_413=1043.333333ns
.PARAM t_a_414=1045ns
.PARAM t_a_415=1048.333333ns
.PARAM t_a_416=1050ns
.PARAM t_a_417=1053.333333ns
.PARAM t_a_418=1055ns
.PARAM t_a_419=1058.333333ns
.PARAM t_a_420=1060ns
.PARAM t_a_421=1063.333333ns
.PARAM t_a_422=1065ns
.PARAM t_a_423=1068.333333ns
.PARAM t_a_424=1070ns
.PARAM t_a_425=1073.333333ns
.PARAM t_a_426=1075ns
.PARAM t_a_427=1078.333333ns
.PARAM t_a_428=1080ns
.PARAM t_a_429=1083.333333ns
.PARAM t_a_430=1085ns
.PARAM t_a_431=1088.333333ns
.PARAM t_a_432=1090ns
.PARAM t_a_433=1093.333333ns
.PARAM t_a_434=1095ns
.PARAM t_a_435=1098.333333ns
.PARAM t_a_436=1100ns
.PARAM t_a_437=1103.333333ns
.PARAM t_a_438=1105ns
.PARAM t_a_439=1108.333333ns
.PARAM t_a_440=1110ns
.PARAM t_a_441=1113.333333ns
.PARAM t_a_442=1115ns
.PARAM t_a_443=1118.333333ns
.PARAM t_a_444=1120ns
.PARAM t_a_445=1123.333333ns
.PARAM t_a_446=1125ns
.PARAM t_a_447=1128.333333ns
.PARAM t_a_448=1130ns
.PARAM t_a_449=1133.333333ns
.PARAM t_a_450=1135ns
.PARAM t_a_451=1138.333333ns
.PARAM t_a_452=1140ns
.PARAM t_a_453=1143.333333ns
.PARAM t_a_454=1145ns
.PARAM t_a_455=1148.333333ns
.PARAM t_a_456=1150ns
.PARAM t_a_457=1153.333333ns
.PARAM t_a_458=1155ns
.PARAM t_a_459=1158.333333ns
.PARAM t_a_460=1160ns
.PARAM t_a_461=1163.333333ns
.PARAM t_a_462=1165ns
.PARAM t_a_463=1168.333333ns
.PARAM t_a_464=1170ns
.PARAM t_a_465=1173.333333ns
.PARAM t_a_466=1175ns
.PARAM t_a_467=1178.333333ns
.PARAM t_a_468=1180ns
.PARAM t_a_469=1183.333333ns
.PARAM t_a_470=1185ns
.PARAM t_a_471=1188.333333ns
.PARAM t_a_472=1190ns
.PARAM t_a_473=1193.333333ns
.PARAM t_a_474=1195ns
.PARAM t_a_475=1198.333333ns
.PARAM t_a_476=1200ns
.PARAM t_a_477=1203.333333ns
.PARAM t_a_478=1205ns
.PARAM t_a_479=1208.333333ns
.PARAM t_a_480=1210ns
.PARAM t_a_481=1213.333333ns
.PARAM t_a_482=1215ns
.PARAM t_a_483=1218.333333ns
.PARAM t_a_484=1220ns
.PARAM t_a_485=1223.333333ns
.PARAM t_a_486=1225ns
.PARAM t_a_487=1228.333333ns
.PARAM t_a_488=1230ns
.PARAM t_a_489=1233.333333ns
.PARAM t_a_490=1235ns
.PARAM t_a_491=1238.333333ns
.PARAM t_a_492=1240ns
.PARAM t_a_493=1243.333333ns
.PARAM t_a_494=1245ns
.PARAM t_a_495=1248.333333ns
.PARAM t_a_496=1250ns
.PARAM t_a_497=1253.333333ns
.PARAM t_a_498=1255ns
.PARAM t_a_499=1258.333333ns
.PARAM t_a_500=1260ns
.PARAM t_a_501=1263.333333ns
.PARAM t_a_502=1265ns
.PARAM t_a_503=1268.333333ns
.PARAM t_a_504=1270ns
.PARAM t_a_505=1273.333333ns
.PARAM t_a_506=1275ns
.PARAM t_a_507=1278.333333ns
.PARAM t_a_508=1280ns
.PARAM t_a_509=1283.333333ns
.PARAM t_a_510=1285ns
.PARAM t_a_511=1288.333333ns
.PARAM t_a_512=1290ns
.PARAM t_a_513=1293.333333ns
.PARAM t_a_514=1295ns
.PARAM t_a_515=1298.333333ns
.PARAM t_a_516=1300ns
.PARAM t_a_517=1303.333333ns
.PARAM t_a_518=1305ns
.PARAM t_a_519=1308.333333ns
.PARAM t_a_520=1310ns
.PARAM t_a_521=1313.333333ns
.PARAM t_a_522=1315ns
.PARAM t_a_523=1318.333333ns
.PARAM t_a_524=1320ns
.PARAM t_a_525=1323.333333ns
.PARAM t_a_526=1325ns
.PARAM t_a_527=1328.333333ns
.PARAM t_a_528=1330ns
.PARAM t_a_529=1333.333333ns
.PARAM t_a_530=1335ns
.PARAM t_a_531=1338.333333ns
.PARAM t_a_532=1340ns
.PARAM t_a_533=1343.333333ns
.PARAM t_a_534=1345ns
.PARAM t_a_535=1348.333333ns
.PARAM t_a_536=1350ns
.PARAM t_a_537=1353.333333ns
.PARAM t_a_538=1355ns
.PARAM t_a_539=1358.333333ns
.PARAM t_a_540=1360ns
.PARAM t_a_541=1363.333333ns
.PARAM t_a_542=1365ns
.PARAM t_a_543=1368.333333ns
.PARAM t_a_544=1370ns
.PARAM t_a_545=1373.333333ns
.PARAM t_a_546=1375ns
.PARAM t_a_547=1378.333333ns
.PARAM t_a_548=1380ns
.PARAM t_a_549=1383.333333ns
.PARAM t_a_550=1385ns
.PARAM t_a_551=1388.333333ns
.PARAM t_a_552=1390ns
.PARAM t_a_553=1393.333333ns
.PARAM t_a_554=1395ns
.PARAM t_a_555=1398.333333ns
.PARAM t_a_556=1400ns
.PARAM t_a_557=1403.333333ns
.PARAM t_a_558=1405ns
.PARAM t_a_559=1408.333333ns
.PARAM t_a_560=1410ns
.PARAM t_a_561=1413.333333ns
.PARAM t_a_562=1415ns
.PARAM t_a_563=1418.333333ns
.PARAM t_a_564=1420ns
.PARAM t_a_565=1423.333333ns
.PARAM t_a_566=1425ns
.PARAM t_a_567=1428.333333ns
.PARAM t_a_568=1430ns
.PARAM t_a_569=1433.333333ns
.PARAM t_a_570=1435ns
.PARAM t_a_571=1438.333333ns
.PARAM t_a_572=1440ns
.PARAM t_a_573=1443.333333ns
.PARAM t_a_574=1445ns
.PARAM t_a_575=1448.333333ns
.PARAM t_a_576=1450ns
.PARAM t_a_577=1453.333333ns
.PARAM t_a_578=1455ns
.PARAM t_a_579=1458.333333ns
.PARAM t_a_580=1460ns
.PARAM t_a_581=1463.333333ns
.PARAM t_a_582=1465ns
.PARAM t_a_583=1468.333333ns
.PARAM t_a_584=1470ns
.PARAM t_a_585=1473.333333ns
.PARAM t_a_586=1475ns
.PARAM t_a_587=1478.333333ns
.PARAM t_a_588=1480ns
.PARAM t_a_589=1483.333333ns
.PARAM t_a_590=1485ns
.PARAM t_a_591=1488.333333ns
.PARAM t_a_592=1490ns
.PARAM t_a_593=1493.333333ns
.PARAM t_a_594=1495ns
.PARAM t_a_595=1498.333333ns
.PARAM t_a_596=1500ns
.PARAM t_a_597=1503.333333ns
.PARAM t_a_598=1505ns
.PARAM t_a_599=1508.333333ns
.PARAM t_a_600=1510ns
.PARAM t_a_601=1513.333333ns
.PARAM t_a_602=1515ns
.PARAM t_a_603=1518.333333ns
.PARAM t_a_604=1520ns
.PARAM t_a_605=1523.333333ns
.PARAM t_a_606=1525ns
.PARAM t_a_607=1528.333333ns
.PARAM t_a_608=1530ns
.PARAM t_a_609=1533.333333ns
.PARAM t_a_610=1535ns
.PARAM t_a_611=1538.333333ns
.PARAM t_a_612=1540ns
.PARAM t_a_613=1543.333333ns
.PARAM t_a_614=1545ns
.PARAM t_a_615=1548.333333ns
.PARAM t_a_616=1550ns
.PARAM t_a_617=1553.333333ns
.PARAM t_a_618=1555ns
.PARAM t_a_619=1558.333333ns
.PARAM t_a_620=1560ns
.PARAM t_a_621=1563.333333ns
.PARAM t_a_622=1565ns
.PARAM t_a_623=1568.333333ns
.PARAM t_a_624=1570ns
.PARAM t_a_625=1573.333333ns
.PARAM t_a_626=1575ns
.PARAM t_a_627=1578.333333ns
.PARAM t_a_628=1580ns
.PARAM t_a_629=1583.333333ns
.PARAM t_a_630=1585ns
.PARAM t_a_631=1588.333333ns
.PARAM t_a_632=1590ns
.PARAM t_a_633=1593.333333ns
.PARAM t_a_634=1595ns
.PARAM t_a_635=1598.333333ns
.PARAM t_a_636=1600ns
.PARAM t_a_637=1603.333333ns
.PARAM t_a_638=1605ns
.PARAM t_a_639=1608.333333ns
.PARAM t_a_640=1610ns
.PARAM t_a_641=1613.333333ns
.PARAM t_a_642=1615ns
.PARAM t_a_643=1618.333333ns
.PARAM t_a_644=1620ns
.PARAM t_a_645=1623.333333ns
.PARAM t_a_646=1625ns
.PARAM t_a_647=1628.333333ns
.PARAM t_a_648=1630ns
.PARAM t_a_649=1633.333333ns
.PARAM t_a_650=1635ns
.PARAM t_a_651=1638.333333ns
.PARAM t_a_652=1640ns
.PARAM t_a_653=1643.333333ns
.PARAM t_a_654=1645ns
.PARAM t_a_655=1648.333333ns
.PARAM t_a_656=1650ns
.PARAM t_a_657=1653.333333ns
.PARAM t_a_658=1655ns
.PARAM t_a_659=1658.333333ns
.PARAM t_a_660=1660ns
.PARAM t_a_661=1663.333333ns
.PARAM t_a_662=1665ns
.PARAM t_a_663=1668.333333ns
.PARAM t_a_664=1670ns
.PARAM t_a_665=1673.333333ns
.PARAM t_a_666=1675ns
.PARAM t_a_667=1678.333333ns
.PARAM t_a_668=1680ns
.PARAM t_a_669=1683.333333ns
.PARAM t_a_670=1685ns
.PARAM t_a_671=1688.333333ns
.PARAM t_a_672=1690ns
.PARAM t_a_673=1693.333333ns
.PARAM t_a_674=1695ns
.PARAM t_a_675=1698.333333ns
.PARAM t_a_676=1700ns
.PARAM t_a_677=1703.333333ns
.PARAM t_a_678=1705ns
.PARAM t_a_679=1708.333333ns
.PARAM t_a_680=1710ns
.PARAM t_a_681=1713.333333ns
.PARAM t_a_682=1715ns
.PARAM t_a_683=1718.333333ns
.PARAM t_a_684=1720ns
.PARAM t_a_685=1723.333333ns
.PARAM t_a_686=1725ns
.PARAM t_a_687=1728.333333ns
.PARAM t_a_688=1730ns
.PARAM t_a_689=1733.333333ns
.PARAM t_a_690=1735ns
.PARAM t_a_691=1738.333333ns
.PARAM t_a_692=1740ns
.PARAM t_a_693=1743.333333ns
.PARAM t_a_694=1745ns
.PARAM t_a_695=1748.333333ns
.PARAM t_a_696=1750ns
.PARAM t_a_697=1753.333333ns
.PARAM t_a_698=1755ns
.PARAM t_a_699=1758.333333ns
.PARAM t_a_700=1760ns
.PARAM t_a_701=1763.333333ns
.PARAM t_a_702=1765ns
.PARAM t_a_703=1768.333333ns
.PARAM t_a_704=1770ns
.PARAM t_a_705=1773.333333ns
.PARAM t_a_706=1775ns
.PARAM t_a_707=1778.333333ns
.PARAM t_a_708=1780ns
.PARAM t_a_709=1783.333333ns
.PARAM t_a_710=1785ns
.PARAM t_a_711=1788.333333ns
.PARAM t_a_712=1790ns
.PARAM t_a_713=1793.333333ns
.PARAM t_a_714=1795ns
.PARAM t_a_715=1798.333333ns
.PARAM t_a_716=1800ns
.PARAM t_a_717=1803.333333ns
.PARAM t_a_718=1805ns
.PARAM t_a_719=1808.333333ns
.PARAM t_a_720=1810ns
.PARAM t_a_721=1813.333333ns
.PARAM t_a_722=1815ns
.PARAM t_a_723=1818.333333ns
.PARAM t_a_724=1820ns
.PARAM t_a_725=1823.333333ns
.PARAM t_a_726=1825ns
.PARAM t_a_727=1828.333333ns
.PARAM t_a_728=1830ns
.PARAM t_a_729=1833.333333ns
.PARAM t_a_730=1835ns
.PARAM t_a_731=1838.333333ns
.PARAM t_a_732=1840ns
.PARAM t_a_733=1843.333333ns
.PARAM t_a_734=1845ns
.PARAM t_a_735=1848.333333ns
.PARAM t_a_736=1850ns
.PARAM t_a_737=1853.333333ns
.PARAM t_a_738=1855ns
.PARAM t_a_739=1858.333333ns
.PARAM t_a_740=1860ns
.PARAM t_a_741=1863.333333ns
.PARAM t_a_742=1865ns
.PARAM t_a_743=1868.333333ns
.PARAM t_a_744=1870ns
.PARAM t_a_745=1873.333333ns
.PARAM t_a_746=1875ns
.PARAM t_a_747=1878.333333ns
.PARAM t_a_748=1880ns
.PARAM t_a_749=1883.333333ns
.PARAM t_a_750=1885ns
.PARAM t_a_751=1888.333333ns
.PARAM t_a_752=1890ns
.PARAM t_a_753=1893.333333ns
.PARAM t_a_754=1895ns
.PARAM t_a_755=1898.333333ns
.PARAM t_a_756=1900ns
.PARAM t_a_757=1903.333333ns
.PARAM t_a_758=1905ns
.PARAM t_a_759=1908.333333ns
.PARAM t_a_760=1910ns
.PARAM t_a_761=1913.333333ns
.PARAM t_a_762=1915ns
.PARAM t_a_763=1918.333333ns
.PARAM t_a_764=1920ns
.PARAM t_a_765=1923.333333ns
.PARAM t_a_766=1925ns
.PARAM t_a_767=1928.333333ns
.PARAM t_a_768=1930ns
.PARAM t_a_769=1933.333333ns
.PARAM t_a_770=1935ns
.PARAM t_a_771=1938.333333ns
.PARAM t_a_772=1940ns
.PARAM t_a_773=1943.333333ns
.PARAM t_a_774=1945ns
.PARAM t_a_775=1948.333333ns
.PARAM t_a_776=1950ns
.PARAM t_a_777=1953.333333ns
.PARAM t_a_778=1955ns
.PARAM t_a_779=1958.333333ns
.PARAM t_a_780=1960ns
.PARAM t_a_781=1963.333333ns
.PARAM t_a_782=1965ns
.PARAM t_a_783=1968.333333ns
.PARAM t_a_784=1970ns
.PARAM t_a_785=1973.333333ns
.PARAM t_a_786=1975ns
.PARAM t_a_787=1978.333333ns
.PARAM t_a_788=1980ns
.PARAM t_a_789=1983.333333ns
.PARAM t_a_790=1985ns
.PARAM t_a_791=1988.333333ns
.PARAM t_a_792=1990ns
.PARAM t_a_793=1993.333333ns
.PARAM t_a_794=1995ns
.PARAM t_a_795=1998.333333ns
.PARAM t_a_796=2000ns
.PARAM t_a_797=2003.333333ns
.PARAM t_a_798=2005ns
.PARAM t_a_799=2008.333333ns
.PARAM t_b_0=9.8ns
.PARAM t_b_1=11.666667ns
.PARAM t_b_2=14.801ns
.PARAM t_b_3=16.666667ns
.PARAM t_b_4=19.802ns
.PARAM t_b_5=21.666667ns
.PARAM t_b_6=24.803ns
.PARAM t_b_7=26.666667ns
.PARAM t_b_8=29.804ns
.PARAM t_b_9=31.666667ns
.PARAM t_b_10=34.805ns
.PARAM t_b_11=36.666667ns
.PARAM t_b_12=39.806ns
.PARAM t_b_13=41.666667ns
.PARAM t_b_14=44.807ns
.PARAM t_b_15=46.666667ns
.PARAM t_b_16=49.808ns
.PARAM t_b_17=51.666667ns
.PARAM t_b_18=54.809ns
.PARAM t_b_19=56.666667ns
.PARAM t_b_20=59.81ns
.PARAM t_b_21=61.666667ns
.PARAM t_b_22=64.811ns
.PARAM t_b_23=66.666667ns
.PARAM t_b_24=69.812ns
.PARAM t_b_25=71.666667ns
.PARAM t_b_26=74.813ns
.PARAM t_b_27=76.666667ns
.PARAM t_b_28=79.814ns
.PARAM t_b_29=81.666667ns
.PARAM t_b_30=84.815ns
.PARAM t_b_31=86.666667ns
.PARAM t_b_32=89.816ns
.PARAM t_b_33=91.666667ns
.PARAM t_b_34=94.817ns
.PARAM t_b_35=96.666667ns
.PARAM t_b_36=99.818ns
.PARAM t_b_37=101.666667ns
.PARAM t_b_38=104.819ns
.PARAM t_b_39=106.666667ns
.PARAM t_b_40=109.82ns
.PARAM t_b_41=111.666667ns
.PARAM t_b_42=114.821ns
.PARAM t_b_43=116.666667ns
.PARAM t_b_44=119.822ns
.PARAM t_b_45=121.666667ns
.PARAM t_b_46=124.823ns
.PARAM t_b_47=126.666667ns
.PARAM t_b_48=129.824ns
.PARAM t_b_49=131.666667ns
.PARAM t_b_50=134.825ns
.PARAM t_b_51=136.666667ns
.PARAM t_b_52=139.826ns
.PARAM t_b_53=141.666667ns
.PARAM t_b_54=144.827ns
.PARAM t_b_55=146.666667ns
.PARAM t_b_56=149.828ns
.PARAM t_b_57=151.666667ns
.PARAM t_b_58=154.829ns
.PARAM t_b_59=156.666667ns
.PARAM t_b_60=159.83ns
.PARAM t_b_61=161.666667ns
.PARAM t_b_62=164.831ns
.PARAM t_b_63=166.666667ns
.PARAM t_b_64=169.832ns
.PARAM t_b_65=171.666667ns
.PARAM t_b_66=174.833ns
.PARAM t_b_67=176.666667ns
.PARAM t_b_68=179.834ns
.PARAM t_b_69=181.666667ns
.PARAM t_b_70=184.835ns
.PARAM t_b_71=186.666667ns
.PARAM t_b_72=189.836ns
.PARAM t_b_73=191.666667ns
.PARAM t_b_74=194.837ns
.PARAM t_b_75=196.666667ns
.PARAM t_b_76=199.838ns
.PARAM t_b_77=201.666667ns
.PARAM t_b_78=204.839ns
.PARAM t_b_79=206.666667ns
.PARAM t_b_80=209.84ns
.PARAM t_b_81=211.666667ns
.PARAM t_b_82=214.841ns
.PARAM t_b_83=216.666667ns
.PARAM t_b_84=219.842ns
.PARAM t_b_85=221.666667ns
.PARAM t_b_86=224.843ns
.PARAM t_b_87=226.666667ns
.PARAM t_b_88=229.844ns
.PARAM t_b_89=231.666667ns
.PARAM t_b_90=234.845ns
.PARAM t_b_91=236.666667ns
.PARAM t_b_92=239.846ns
.PARAM t_b_93=241.666667ns
.PARAM t_b_94=244.847ns
.PARAM t_b_95=246.666667ns
.PARAM t_b_96=249.848ns
.PARAM t_b_97=251.666667ns
.PARAM t_b_98=254.849ns
.PARAM t_b_99=256.666667ns
.PARAM t_b_100=259.85ns
.PARAM t_b_101=261.666667ns
.PARAM t_b_102=264.851ns
.PARAM t_b_103=266.666667ns
.PARAM t_b_104=269.852ns
.PARAM t_b_105=271.666667ns
.PARAM t_b_106=274.853ns
.PARAM t_b_107=276.666667ns
.PARAM t_b_108=279.854ns
.PARAM t_b_109=281.666667ns
.PARAM t_b_110=284.855ns
.PARAM t_b_111=286.666667ns
.PARAM t_b_112=289.856ns
.PARAM t_b_113=291.666667ns
.PARAM t_b_114=294.857ns
.PARAM t_b_115=296.666667ns
.PARAM t_b_116=299.858ns
.PARAM t_b_117=301.666667ns
.PARAM t_b_118=304.859ns
.PARAM t_b_119=306.666667ns
.PARAM t_b_120=309.86ns
.PARAM t_b_121=311.666667ns
.PARAM t_b_122=314.861ns
.PARAM t_b_123=316.666667ns
.PARAM t_b_124=319.862ns
.PARAM t_b_125=321.666667ns
.PARAM t_b_126=324.863ns
.PARAM t_b_127=326.666667ns
.PARAM t_b_128=329.864ns
.PARAM t_b_129=331.666667ns
.PARAM t_b_130=334.865ns
.PARAM t_b_131=336.666667ns
.PARAM t_b_132=339.866ns
.PARAM t_b_133=341.666667ns
.PARAM t_b_134=344.867ns
.PARAM t_b_135=346.666667ns
.PARAM t_b_136=349.868ns
.PARAM t_b_137=351.666667ns
.PARAM t_b_138=354.869ns
.PARAM t_b_139=356.666667ns
.PARAM t_b_140=359.87ns
.PARAM t_b_141=361.666667ns
.PARAM t_b_142=364.871ns
.PARAM t_b_143=366.666667ns
.PARAM t_b_144=369.872ns
.PARAM t_b_145=371.666667ns
.PARAM t_b_146=374.873ns
.PARAM t_b_147=376.666667ns
.PARAM t_b_148=379.874ns
.PARAM t_b_149=381.666667ns
.PARAM t_b_150=384.875ns
.PARAM t_b_151=386.666667ns
.PARAM t_b_152=389.876ns
.PARAM t_b_153=391.666667ns
.PARAM t_b_154=394.877ns
.PARAM t_b_155=396.666667ns
.PARAM t_b_156=399.878ns
.PARAM t_b_157=401.666667ns
.PARAM t_b_158=404.879ns
.PARAM t_b_159=406.666667ns
.PARAM t_b_160=409.88ns
.PARAM t_b_161=411.666667ns
.PARAM t_b_162=414.881ns
.PARAM t_b_163=416.666667ns
.PARAM t_b_164=419.882ns
.PARAM t_b_165=421.666667ns
.PARAM t_b_166=424.883ns
.PARAM t_b_167=426.666667ns
.PARAM t_b_168=429.884ns
.PARAM t_b_169=431.666667ns
.PARAM t_b_170=434.885ns
.PARAM t_b_171=436.666667ns
.PARAM t_b_172=439.886ns
.PARAM t_b_173=441.666667ns
.PARAM t_b_174=444.887ns
.PARAM t_b_175=446.666667ns
.PARAM t_b_176=449.888ns
.PARAM t_b_177=451.666667ns
.PARAM t_b_178=454.889ns
.PARAM t_b_179=456.666667ns
.PARAM t_b_180=459.89ns
.PARAM t_b_181=461.666667ns
.PARAM t_b_182=464.891ns
.PARAM t_b_183=466.666667ns
.PARAM t_b_184=469.892ns
.PARAM t_b_185=471.666667ns
.PARAM t_b_186=474.893ns
.PARAM t_b_187=476.666667ns
.PARAM t_b_188=479.894ns
.PARAM t_b_189=481.666667ns
.PARAM t_b_190=484.895ns
.PARAM t_b_191=486.666667ns
.PARAM t_b_192=489.896ns
.PARAM t_b_193=491.666667ns
.PARAM t_b_194=494.897ns
.PARAM t_b_195=496.666667ns
.PARAM t_b_196=499.898ns
.PARAM t_b_197=501.666667ns
.PARAM t_b_198=504.899ns
.PARAM t_b_199=506.666667ns
.PARAM t_b_200=509.9ns
.PARAM t_b_201=511.666667ns
.PARAM t_b_202=514.901ns
.PARAM t_b_203=516.666667ns
.PARAM t_b_204=519.902ns
.PARAM t_b_205=521.666667ns
.PARAM t_b_206=524.903ns
.PARAM t_b_207=526.666667ns
.PARAM t_b_208=529.904ns
.PARAM t_b_209=531.666667ns
.PARAM t_b_210=534.905ns
.PARAM t_b_211=536.666667ns
.PARAM t_b_212=539.906ns
.PARAM t_b_213=541.666667ns
.PARAM t_b_214=544.907ns
.PARAM t_b_215=546.666667ns
.PARAM t_b_216=549.908ns
.PARAM t_b_217=551.666667ns
.PARAM t_b_218=554.909ns
.PARAM t_b_219=556.666667ns
.PARAM t_b_220=559.91ns
.PARAM t_b_221=561.666667ns
.PARAM t_b_222=564.911ns
.PARAM t_b_223=566.666667ns
.PARAM t_b_224=569.912ns
.PARAM t_b_225=571.666667ns
.PARAM t_b_226=574.913ns
.PARAM t_b_227=576.666667ns
.PARAM t_b_228=579.914ns
.PARAM t_b_229=581.666667ns
.PARAM t_b_230=584.915ns
.PARAM t_b_231=586.666667ns
.PARAM t_b_232=589.916ns
.PARAM t_b_233=591.666667ns
.PARAM t_b_234=594.917ns
.PARAM t_b_235=596.666667ns
.PARAM t_b_236=599.918ns
.PARAM t_b_237=601.666667ns
.PARAM t_b_238=604.919ns
.PARAM t_b_239=606.666667ns
.PARAM t_b_240=609.92ns
.PARAM t_b_241=611.666667ns
.PARAM t_b_242=614.921ns
.PARAM t_b_243=616.666667ns
.PARAM t_b_244=619.922ns
.PARAM t_b_245=621.666667ns
.PARAM t_b_246=624.923ns
.PARAM t_b_247=626.666667ns
.PARAM t_b_248=629.924ns
.PARAM t_b_249=631.666667ns
.PARAM t_b_250=634.925ns
.PARAM t_b_251=636.666667ns
.PARAM t_b_252=639.926ns
.PARAM t_b_253=641.666667ns
.PARAM t_b_254=644.927ns
.PARAM t_b_255=646.666667ns
.PARAM t_b_256=649.928ns
.PARAM t_b_257=651.666667ns
.PARAM t_b_258=654.929ns
.PARAM t_b_259=656.666667ns
.PARAM t_b_260=659.93ns
.PARAM t_b_261=661.666667ns
.PARAM t_b_262=664.931ns
.PARAM t_b_263=666.666667ns
.PARAM t_b_264=669.932ns
.PARAM t_b_265=671.666667ns
.PARAM t_b_266=674.933ns
.PARAM t_b_267=676.666667ns
.PARAM t_b_268=679.934ns
.PARAM t_b_269=681.666667ns
.PARAM t_b_270=684.935ns
.PARAM t_b_271=686.666667ns
.PARAM t_b_272=689.936ns
.PARAM t_b_273=691.666667ns
.PARAM t_b_274=694.937ns
.PARAM t_b_275=696.666667ns
.PARAM t_b_276=699.938ns
.PARAM t_b_277=701.666667ns
.PARAM t_b_278=704.939ns
.PARAM t_b_279=706.666667ns
.PARAM t_b_280=709.94ns
.PARAM t_b_281=711.666667ns
.PARAM t_b_282=714.941ns
.PARAM t_b_283=716.666667ns
.PARAM t_b_284=719.942ns
.PARAM t_b_285=721.666667ns
.PARAM t_b_286=724.943ns
.PARAM t_b_287=726.666667ns
.PARAM t_b_288=729.944ns
.PARAM t_b_289=731.666667ns
.PARAM t_b_290=734.945ns
.PARAM t_b_291=736.666667ns
.PARAM t_b_292=739.946ns
.PARAM t_b_293=741.666667ns
.PARAM t_b_294=744.947ns
.PARAM t_b_295=746.666667ns
.PARAM t_b_296=749.948ns
.PARAM t_b_297=751.666667ns
.PARAM t_b_298=754.949ns
.PARAM t_b_299=756.666667ns
.PARAM t_b_300=759.95ns
.PARAM t_b_301=761.666667ns
.PARAM t_b_302=764.951ns
.PARAM t_b_303=766.666667ns
.PARAM t_b_304=769.952ns
.PARAM t_b_305=771.666667ns
.PARAM t_b_306=774.953ns
.PARAM t_b_307=776.666667ns
.PARAM t_b_308=779.954ns
.PARAM t_b_309=781.666667ns
.PARAM t_b_310=784.955ns
.PARAM t_b_311=786.666667ns
.PARAM t_b_312=789.956ns
.PARAM t_b_313=791.666667ns
.PARAM t_b_314=794.957ns
.PARAM t_b_315=796.666667ns
.PARAM t_b_316=799.958ns
.PARAM t_b_317=801.666667ns
.PARAM t_b_318=804.959ns
.PARAM t_b_319=806.666667ns
.PARAM t_b_320=809.96ns
.PARAM t_b_321=811.666667ns
.PARAM t_b_322=814.961ns
.PARAM t_b_323=816.666667ns
.PARAM t_b_324=819.962ns
.PARAM t_b_325=821.666667ns
.PARAM t_b_326=824.963ns
.PARAM t_b_327=826.666667ns
.PARAM t_b_328=829.964ns
.PARAM t_b_329=831.666667ns
.PARAM t_b_330=834.965ns
.PARAM t_b_331=836.666667ns
.PARAM t_b_332=839.966ns
.PARAM t_b_333=841.666667ns
.PARAM t_b_334=844.967ns
.PARAM t_b_335=846.666667ns
.PARAM t_b_336=849.968ns
.PARAM t_b_337=851.666667ns
.PARAM t_b_338=854.969ns
.PARAM t_b_339=856.666667ns
.PARAM t_b_340=859.97ns
.PARAM t_b_341=861.666667ns
.PARAM t_b_342=864.971ns
.PARAM t_b_343=866.666667ns
.PARAM t_b_344=869.972ns
.PARAM t_b_345=871.666667ns
.PARAM t_b_346=874.973ns
.PARAM t_b_347=876.666667ns
.PARAM t_b_348=879.974ns
.PARAM t_b_349=881.666667ns
.PARAM t_b_350=884.975ns
.PARAM t_b_351=886.666667ns
.PARAM t_b_352=889.976ns
.PARAM t_b_353=891.666667ns
.PARAM t_b_354=894.977ns
.PARAM t_b_355=896.666667ns
.PARAM t_b_356=899.978ns
.PARAM t_b_357=901.666667ns
.PARAM t_b_358=904.979ns
.PARAM t_b_359=906.666667ns
.PARAM t_b_360=909.98ns
.PARAM t_b_361=911.666667ns
.PARAM t_b_362=914.981ns
.PARAM t_b_363=916.666667ns
.PARAM t_b_364=919.982ns
.PARAM t_b_365=921.666667ns
.PARAM t_b_366=924.983ns
.PARAM t_b_367=926.666667ns
.PARAM t_b_368=929.984ns
.PARAM t_b_369=931.666667ns
.PARAM t_b_370=934.985ns
.PARAM t_b_371=936.666667ns
.PARAM t_b_372=939.986ns
.PARAM t_b_373=941.666667ns
.PARAM t_b_374=944.987ns
.PARAM t_b_375=946.666667ns
.PARAM t_b_376=949.988ns
.PARAM t_b_377=951.666667ns
.PARAM t_b_378=954.989ns
.PARAM t_b_379=956.666667ns
.PARAM t_b_380=959.99ns
.PARAM t_b_381=961.666667ns
.PARAM t_b_382=964.991ns
.PARAM t_b_383=966.666667ns
.PARAM t_b_384=969.992ns
.PARAM t_b_385=971.666667ns
.PARAM t_b_386=974.993ns
.PARAM t_b_387=976.666667ns
.PARAM t_b_388=979.994ns
.PARAM t_b_389=981.666667ns
.PARAM t_b_390=984.995ns
.PARAM t_b_391=986.666667ns
.PARAM t_b_392=989.996ns
.PARAM t_b_393=991.666667ns
.PARAM t_b_394=994.997ns
.PARAM t_b_395=996.666667ns
.PARAM t_b_396=999.998ns
.PARAM t_b_397=1001.666667ns
.PARAM t_b_398=1004.999ns
.PARAM t_b_399=1006.666667ns
.PARAM t_b_400=1010.0ns
.PARAM t_b_401=1011.666667ns
.PARAM t_b_402=1015.001ns
.PARAM t_b_403=1016.666667ns
.PARAM t_b_404=1020.002ns
.PARAM t_b_405=1021.666667ns
.PARAM t_b_406=1025.003ns
.PARAM t_b_407=1026.666667ns
.PARAM t_b_408=1030.004ns
.PARAM t_b_409=1031.666667ns
.PARAM t_b_410=1035.005ns
.PARAM t_b_411=1036.666667ns
.PARAM t_b_412=1040.006ns
.PARAM t_b_413=1041.666667ns
.PARAM t_b_414=1045.007ns
.PARAM t_b_415=1046.666667ns
.PARAM t_b_416=1050.008ns
.PARAM t_b_417=1051.666667ns
.PARAM t_b_418=1055.009ns
.PARAM t_b_419=1056.666667ns
.PARAM t_b_420=1060.01ns
.PARAM t_b_421=1061.666667ns
.PARAM t_b_422=1065.011ns
.PARAM t_b_423=1066.666667ns
.PARAM t_b_424=1070.012ns
.PARAM t_b_425=1071.666667ns
.PARAM t_b_426=1075.013ns
.PARAM t_b_427=1076.666667ns
.PARAM t_b_428=1080.014ns
.PARAM t_b_429=1081.666667ns
.PARAM t_b_430=1085.015ns
.PARAM t_b_431=1086.666667ns
.PARAM t_b_432=1090.016ns
.PARAM t_b_433=1091.666667ns
.PARAM t_b_434=1095.017ns
.PARAM t_b_435=1096.666667ns
.PARAM t_b_436=1100.018ns
.PARAM t_b_437=1101.666667ns
.PARAM t_b_438=1105.019ns
.PARAM t_b_439=1106.666667ns
.PARAM t_b_440=1110.02ns
.PARAM t_b_441=1111.666667ns
.PARAM t_b_442=1115.021ns
.PARAM t_b_443=1116.666667ns
.PARAM t_b_444=1120.022ns
.PARAM t_b_445=1121.666667ns
.PARAM t_b_446=1125.023ns
.PARAM t_b_447=1126.666667ns
.PARAM t_b_448=1130.024ns
.PARAM t_b_449=1131.666667ns
.PARAM t_b_450=1135.025ns
.PARAM t_b_451=1136.666667ns
.PARAM t_b_452=1140.026ns
.PARAM t_b_453=1141.666667ns
.PARAM t_b_454=1145.027ns
.PARAM t_b_455=1146.666667ns
.PARAM t_b_456=1150.028ns
.PARAM t_b_457=1151.666667ns
.PARAM t_b_458=1155.029ns
.PARAM t_b_459=1156.666667ns
.PARAM t_b_460=1160.03ns
.PARAM t_b_461=1161.666667ns
.PARAM t_b_462=1165.031ns
.PARAM t_b_463=1166.666667ns
.PARAM t_b_464=1170.032ns
.PARAM t_b_465=1171.666667ns
.PARAM t_b_466=1175.033ns
.PARAM t_b_467=1176.666667ns
.PARAM t_b_468=1180.034ns
.PARAM t_b_469=1181.666667ns
.PARAM t_b_470=1185.035ns
.PARAM t_b_471=1186.666667ns
.PARAM t_b_472=1190.036ns
.PARAM t_b_473=1191.666667ns
.PARAM t_b_474=1195.037ns
.PARAM t_b_475=1196.666667ns
.PARAM t_b_476=1200.038ns
.PARAM t_b_477=1201.666667ns
.PARAM t_b_478=1205.039ns
.PARAM t_b_479=1206.666667ns
.PARAM t_b_480=1210.04ns
.PARAM t_b_481=1211.666667ns
.PARAM t_b_482=1215.041ns
.PARAM t_b_483=1216.666667ns
.PARAM t_b_484=1220.042ns
.PARAM t_b_485=1221.666667ns
.PARAM t_b_486=1225.043ns
.PARAM t_b_487=1226.666667ns
.PARAM t_b_488=1230.044ns
.PARAM t_b_489=1231.666667ns
.PARAM t_b_490=1235.045ns
.PARAM t_b_491=1236.666667ns
.PARAM t_b_492=1240.046ns
.PARAM t_b_493=1241.666667ns
.PARAM t_b_494=1245.047ns
.PARAM t_b_495=1246.666667ns
.PARAM t_b_496=1250.048ns
.PARAM t_b_497=1251.666667ns
.PARAM t_b_498=1255.049ns
.PARAM t_b_499=1256.666667ns
.PARAM t_b_500=1260.05ns
.PARAM t_b_501=1261.666667ns
.PARAM t_b_502=1265.051ns
.PARAM t_b_503=1266.666667ns
.PARAM t_b_504=1270.052ns
.PARAM t_b_505=1271.666667ns
.PARAM t_b_506=1275.053ns
.PARAM t_b_507=1276.666667ns
.PARAM t_b_508=1280.054ns
.PARAM t_b_509=1281.666667ns
.PARAM t_b_510=1285.055ns
.PARAM t_b_511=1286.666667ns
.PARAM t_b_512=1290.056ns
.PARAM t_b_513=1291.666667ns
.PARAM t_b_514=1295.057ns
.PARAM t_b_515=1296.666667ns
.PARAM t_b_516=1300.058ns
.PARAM t_b_517=1301.666667ns
.PARAM t_b_518=1305.059ns
.PARAM t_b_519=1306.666667ns
.PARAM t_b_520=1310.06ns
.PARAM t_b_521=1311.666667ns
.PARAM t_b_522=1315.061ns
.PARAM t_b_523=1316.666667ns
.PARAM t_b_524=1320.062ns
.PARAM t_b_525=1321.666667ns
.PARAM t_b_526=1325.063ns
.PARAM t_b_527=1326.666667ns
.PARAM t_b_528=1330.064ns
.PARAM t_b_529=1331.666667ns
.PARAM t_b_530=1335.065ns
.PARAM t_b_531=1336.666667ns
.PARAM t_b_532=1340.066ns
.PARAM t_b_533=1341.666667ns
.PARAM t_b_534=1345.067ns
.PARAM t_b_535=1346.666667ns
.PARAM t_b_536=1350.068ns
.PARAM t_b_537=1351.666667ns
.PARAM t_b_538=1355.069ns
.PARAM t_b_539=1356.666667ns
.PARAM t_b_540=1360.07ns
.PARAM t_b_541=1361.666667ns
.PARAM t_b_542=1365.071ns
.PARAM t_b_543=1366.666667ns
.PARAM t_b_544=1370.072ns
.PARAM t_b_545=1371.666667ns
.PARAM t_b_546=1375.073ns
.PARAM t_b_547=1376.666667ns
.PARAM t_b_548=1380.074ns
.PARAM t_b_549=1381.666667ns
.PARAM t_b_550=1385.075ns
.PARAM t_b_551=1386.666667ns
.PARAM t_b_552=1390.076ns
.PARAM t_b_553=1391.666667ns
.PARAM t_b_554=1395.077ns
.PARAM t_b_555=1396.666667ns
.PARAM t_b_556=1400.078ns
.PARAM t_b_557=1401.666667ns
.PARAM t_b_558=1405.079ns
.PARAM t_b_559=1406.666667ns
.PARAM t_b_560=1410.08ns
.PARAM t_b_561=1411.666667ns
.PARAM t_b_562=1415.081ns
.PARAM t_b_563=1416.666667ns
.PARAM t_b_564=1420.082ns
.PARAM t_b_565=1421.666667ns
.PARAM t_b_566=1425.083ns
.PARAM t_b_567=1426.666667ns
.PARAM t_b_568=1430.084ns
.PARAM t_b_569=1431.666667ns
.PARAM t_b_570=1435.085ns
.PARAM t_b_571=1436.666667ns
.PARAM t_b_572=1440.086ns
.PARAM t_b_573=1441.666667ns
.PARAM t_b_574=1445.087ns
.PARAM t_b_575=1446.666667ns
.PARAM t_b_576=1450.088ns
.PARAM t_b_577=1451.666667ns
.PARAM t_b_578=1455.089ns
.PARAM t_b_579=1456.666667ns
.PARAM t_b_580=1460.09ns
.PARAM t_b_581=1461.666667ns
.PARAM t_b_582=1465.091ns
.PARAM t_b_583=1466.666667ns
.PARAM t_b_584=1470.092ns
.PARAM t_b_585=1471.666667ns
.PARAM t_b_586=1475.093ns
.PARAM t_b_587=1476.666667ns
.PARAM t_b_588=1480.094ns
.PARAM t_b_589=1481.666667ns
.PARAM t_b_590=1485.095ns
.PARAM t_b_591=1486.666667ns
.PARAM t_b_592=1490.096ns
.PARAM t_b_593=1491.666667ns
.PARAM t_b_594=1495.097ns
.PARAM t_b_595=1496.666667ns
.PARAM t_b_596=1500.098ns
.PARAM t_b_597=1501.666667ns
.PARAM t_b_598=1505.099ns
.PARAM t_b_599=1506.666667ns
.PARAM t_b_600=1510.1ns
.PARAM t_b_601=1511.666667ns
.PARAM t_b_602=1515.101ns
.PARAM t_b_603=1516.666667ns
.PARAM t_b_604=1520.102ns
.PARAM t_b_605=1521.666667ns
.PARAM t_b_606=1525.103ns
.PARAM t_b_607=1526.666667ns
.PARAM t_b_608=1530.104ns
.PARAM t_b_609=1531.666667ns
.PARAM t_b_610=1535.105ns
.PARAM t_b_611=1536.666667ns
.PARAM t_b_612=1540.106ns
.PARAM t_b_613=1541.666667ns
.PARAM t_b_614=1545.107ns
.PARAM t_b_615=1546.666667ns
.PARAM t_b_616=1550.108ns
.PARAM t_b_617=1551.666667ns
.PARAM t_b_618=1555.109ns
.PARAM t_b_619=1556.666667ns
.PARAM t_b_620=1560.11ns
.PARAM t_b_621=1561.666667ns
.PARAM t_b_622=1565.111ns
.PARAM t_b_623=1566.666667ns
.PARAM t_b_624=1570.112ns
.PARAM t_b_625=1571.666667ns
.PARAM t_b_626=1575.113ns
.PARAM t_b_627=1576.666667ns
.PARAM t_b_628=1580.114ns
.PARAM t_b_629=1581.666667ns
.PARAM t_b_630=1585.115ns
.PARAM t_b_631=1586.666667ns
.PARAM t_b_632=1590.116ns
.PARAM t_b_633=1591.666667ns
.PARAM t_b_634=1595.117ns
.PARAM t_b_635=1596.666667ns
.PARAM t_b_636=1600.118ns
.PARAM t_b_637=1601.666667ns
.PARAM t_b_638=1605.119ns
.PARAM t_b_639=1606.666667ns
.PARAM t_b_640=1610.12ns
.PARAM t_b_641=1611.666667ns
.PARAM t_b_642=1615.121ns
.PARAM t_b_643=1616.666667ns
.PARAM t_b_644=1620.122ns
.PARAM t_b_645=1621.666667ns
.PARAM t_b_646=1625.123ns
.PARAM t_b_647=1626.666667ns
.PARAM t_b_648=1630.124ns
.PARAM t_b_649=1631.666667ns
.PARAM t_b_650=1635.125ns
.PARAM t_b_651=1636.666667ns
.PARAM t_b_652=1640.126ns
.PARAM t_b_653=1641.666667ns
.PARAM t_b_654=1645.127ns
.PARAM t_b_655=1646.666667ns
.PARAM t_b_656=1650.128ns
.PARAM t_b_657=1651.666667ns
.PARAM t_b_658=1655.129ns
.PARAM t_b_659=1656.666667ns
.PARAM t_b_660=1660.13ns
.PARAM t_b_661=1661.666667ns
.PARAM t_b_662=1665.131ns
.PARAM t_b_663=1666.666667ns
.PARAM t_b_664=1670.132ns
.PARAM t_b_665=1671.666667ns
.PARAM t_b_666=1675.133ns
.PARAM t_b_667=1676.666667ns
.PARAM t_b_668=1680.134ns
.PARAM t_b_669=1681.666667ns
.PARAM t_b_670=1685.135ns
.PARAM t_b_671=1686.666667ns
.PARAM t_b_672=1690.136ns
.PARAM t_b_673=1691.666667ns
.PARAM t_b_674=1695.137ns
.PARAM t_b_675=1696.666667ns
.PARAM t_b_676=1700.138ns
.PARAM t_b_677=1701.666667ns
.PARAM t_b_678=1705.139ns
.PARAM t_b_679=1706.666667ns
.PARAM t_b_680=1710.14ns
.PARAM t_b_681=1711.666667ns
.PARAM t_b_682=1715.141ns
.PARAM t_b_683=1716.666667ns
.PARAM t_b_684=1720.142ns
.PARAM t_b_685=1721.666667ns
.PARAM t_b_686=1725.143ns
.PARAM t_b_687=1726.666667ns
.PARAM t_b_688=1730.144ns
.PARAM t_b_689=1731.666667ns
.PARAM t_b_690=1735.145ns
.PARAM t_b_691=1736.666667ns
.PARAM t_b_692=1740.146ns
.PARAM t_b_693=1741.666667ns
.PARAM t_b_694=1745.147ns
.PARAM t_b_695=1746.666667ns
.PARAM t_b_696=1750.148ns
.PARAM t_b_697=1751.666667ns
.PARAM t_b_698=1755.149ns
.PARAM t_b_699=1756.666667ns
.PARAM t_b_700=1760.15ns
.PARAM t_b_701=1761.666667ns
.PARAM t_b_702=1765.151ns
.PARAM t_b_703=1766.666667ns
.PARAM t_b_704=1770.152ns
.PARAM t_b_705=1771.666667ns
.PARAM t_b_706=1775.153ns
.PARAM t_b_707=1776.666667ns
.PARAM t_b_708=1780.154ns
.PARAM t_b_709=1781.666667ns
.PARAM t_b_710=1785.155ns
.PARAM t_b_711=1786.666667ns
.PARAM t_b_712=1790.156ns
.PARAM t_b_713=1791.666667ns
.PARAM t_b_714=1795.157ns
.PARAM t_b_715=1796.666667ns
.PARAM t_b_716=1800.158ns
.PARAM t_b_717=1801.666667ns
.PARAM t_b_718=1805.159ns
.PARAM t_b_719=1806.666667ns
.PARAM t_b_720=1810.16ns
.PARAM t_b_721=1811.666667ns
.PARAM t_b_722=1815.161ns
.PARAM t_b_723=1816.666667ns
.PARAM t_b_724=1820.162ns
.PARAM t_b_725=1821.666667ns
.PARAM t_b_726=1825.163ns
.PARAM t_b_727=1826.666667ns
.PARAM t_b_728=1830.164ns
.PARAM t_b_729=1831.666667ns
.PARAM t_b_730=1835.165ns
.PARAM t_b_731=1836.666667ns
.PARAM t_b_732=1840.166ns
.PARAM t_b_733=1841.666667ns
.PARAM t_b_734=1845.167ns
.PARAM t_b_735=1846.666667ns
.PARAM t_b_736=1850.168ns
.PARAM t_b_737=1851.666667ns
.PARAM t_b_738=1855.169ns
.PARAM t_b_739=1856.666667ns
.PARAM t_b_740=1860.17ns
.PARAM t_b_741=1861.666667ns
.PARAM t_b_742=1865.171ns
.PARAM t_b_743=1866.666667ns
.PARAM t_b_744=1870.172ns
.PARAM t_b_745=1871.666667ns
.PARAM t_b_746=1875.173ns
.PARAM t_b_747=1876.666667ns
.PARAM t_b_748=1880.174ns
.PARAM t_b_749=1881.666667ns
.PARAM t_b_750=1885.175ns
.PARAM t_b_751=1886.666667ns
.PARAM t_b_752=1890.176ns
.PARAM t_b_753=1891.666667ns
.PARAM t_b_754=1895.177ns
.PARAM t_b_755=1896.666667ns
.PARAM t_b_756=1900.178ns
.PARAM t_b_757=1901.666667ns
.PARAM t_b_758=1905.179ns
.PARAM t_b_759=1906.666667ns
.PARAM t_b_760=1910.18ns
.PARAM t_b_761=1911.666667ns
.PARAM t_b_762=1915.181ns
.PARAM t_b_763=1916.666667ns
.PARAM t_b_764=1920.182ns
.PARAM t_b_765=1921.666667ns
.PARAM t_b_766=1925.183ns
.PARAM t_b_767=1926.666667ns
.PARAM t_b_768=1930.184ns
.PARAM t_b_769=1931.666667ns
.PARAM t_b_770=1935.185ns
.PARAM t_b_771=1936.666667ns
.PARAM t_b_772=1940.186ns
.PARAM t_b_773=1941.666667ns
.PARAM t_b_774=1945.187ns
.PARAM t_b_775=1946.666667ns
.PARAM t_b_776=1950.188ns
.PARAM t_b_777=1951.666667ns
.PARAM t_b_778=1955.189ns
.PARAM t_b_779=1956.666667ns
.PARAM t_b_780=1960.19ns
.PARAM t_b_781=1961.666667ns
.PARAM t_b_782=1965.191ns
.PARAM t_b_783=1966.666667ns
.PARAM t_b_784=1970.192ns
.PARAM t_b_785=1971.666667ns
.PARAM t_b_786=1975.193ns
.PARAM t_b_787=1976.666667ns
.PARAM t_b_788=1980.194ns
.PARAM t_b_789=1981.666667ns
.PARAM t_b_790=1985.195ns
.PARAM t_b_791=1986.666667ns
.PARAM t_b_792=1990.196ns
.PARAM t_b_793=1991.666667ns
.PARAM t_b_794=1995.197ns
.PARAM t_b_795=1996.666667ns
.PARAM t_b_796=2000.198ns
.PARAM t_b_797=2001.666667ns
.PARAM t_b_798=2005.199ns
.PARAM t_b_799=2006.666667ns



VINA Input_A GND PWL 0ns baseVal t_init0 baseVal 't_init0+slope' peakVal t_init1 peakVal 't_init1+slope' baseVal
+ t_a_0 baseVal 't_a_0+slope' peakVal
+ t_a_1 peakVal 't_a_1+slope' baseVal
+ t_a_2 baseVal 't_a_2+slope' peakVal
+ t_a_3 peakVal 't_a_3+slope' baseVal
+ t_a_4 baseVal 't_a_4+slope' peakVal
+ t_a_5 peakVal 't_a_5+slope' baseVal
+ t_a_6 baseVal 't_a_6+slope' peakVal
+ t_a_7 peakVal 't_a_7+slope' baseVal
+ t_a_8 baseVal 't_a_8+slope' peakVal
+ t_a_9 peakVal 't_a_9+slope' baseVal
+ t_a_10 baseVal 't_a_10+slope' peakVal
+ t_a_11 peakVal 't_a_11+slope' baseVal
+ t_a_12 baseVal 't_a_12+slope' peakVal
+ t_a_13 peakVal 't_a_13+slope' baseVal
+ t_a_14 baseVal 't_a_14+slope' peakVal
+ t_a_15 peakVal 't_a_15+slope' baseVal
+ t_a_16 baseVal 't_a_16+slope' peakVal
+ t_a_17 peakVal 't_a_17+slope' baseVal
+ t_a_18 baseVal 't_a_18+slope' peakVal
+ t_a_19 peakVal 't_a_19+slope' baseVal
+ t_a_20 baseVal 't_a_20+slope' peakVal
+ t_a_21 peakVal 't_a_21+slope' baseVal
+ t_a_22 baseVal 't_a_22+slope' peakVal
+ t_a_23 peakVal 't_a_23+slope' baseVal
+ t_a_24 baseVal 't_a_24+slope' peakVal
+ t_a_25 peakVal 't_a_25+slope' baseVal
+ t_a_26 baseVal 't_a_26+slope' peakVal
+ t_a_27 peakVal 't_a_27+slope' baseVal
+ t_a_28 baseVal 't_a_28+slope' peakVal
+ t_a_29 peakVal 't_a_29+slope' baseVal
+ t_a_30 baseVal 't_a_30+slope' peakVal
+ t_a_31 peakVal 't_a_31+slope' baseVal
+ t_a_32 baseVal 't_a_32+slope' peakVal
+ t_a_33 peakVal 't_a_33+slope' baseVal
+ t_a_34 baseVal 't_a_34+slope' peakVal
+ t_a_35 peakVal 't_a_35+slope' baseVal
+ t_a_36 baseVal 't_a_36+slope' peakVal
+ t_a_37 peakVal 't_a_37+slope' baseVal
+ t_a_38 baseVal 't_a_38+slope' peakVal
+ t_a_39 peakVal 't_a_39+slope' baseVal
+ t_a_40 baseVal 't_a_40+slope' peakVal
+ t_a_41 peakVal 't_a_41+slope' baseVal
+ t_a_42 baseVal 't_a_42+slope' peakVal
+ t_a_43 peakVal 't_a_43+slope' baseVal
+ t_a_44 baseVal 't_a_44+slope' peakVal
+ t_a_45 peakVal 't_a_45+slope' baseVal
+ t_a_46 baseVal 't_a_46+slope' peakVal
+ t_a_47 peakVal 't_a_47+slope' baseVal
+ t_a_48 baseVal 't_a_48+slope' peakVal
+ t_a_49 peakVal 't_a_49+slope' baseVal
+ t_a_50 baseVal 't_a_50+slope' peakVal
+ t_a_51 peakVal 't_a_51+slope' baseVal
+ t_a_52 baseVal 't_a_52+slope' peakVal
+ t_a_53 peakVal 't_a_53+slope' baseVal
+ t_a_54 baseVal 't_a_54+slope' peakVal
+ t_a_55 peakVal 't_a_55+slope' baseVal
+ t_a_56 baseVal 't_a_56+slope' peakVal
+ t_a_57 peakVal 't_a_57+slope' baseVal
+ t_a_58 baseVal 't_a_58+slope' peakVal
+ t_a_59 peakVal 't_a_59+slope' baseVal
+ t_a_60 baseVal 't_a_60+slope' peakVal
+ t_a_61 peakVal 't_a_61+slope' baseVal
+ t_a_62 baseVal 't_a_62+slope' peakVal
+ t_a_63 peakVal 't_a_63+slope' baseVal
+ t_a_64 baseVal 't_a_64+slope' peakVal
+ t_a_65 peakVal 't_a_65+slope' baseVal
+ t_a_66 baseVal 't_a_66+slope' peakVal
+ t_a_67 peakVal 't_a_67+slope' baseVal
+ t_a_68 baseVal 't_a_68+slope' peakVal
+ t_a_69 peakVal 't_a_69+slope' baseVal
+ t_a_70 baseVal 't_a_70+slope' peakVal
+ t_a_71 peakVal 't_a_71+slope' baseVal
+ t_a_72 baseVal 't_a_72+slope' peakVal
+ t_a_73 peakVal 't_a_73+slope' baseVal
+ t_a_74 baseVal 't_a_74+slope' peakVal
+ t_a_75 peakVal 't_a_75+slope' baseVal
+ t_a_76 baseVal 't_a_76+slope' peakVal
+ t_a_77 peakVal 't_a_77+slope' baseVal
+ t_a_78 baseVal 't_a_78+slope' peakVal
+ t_a_79 peakVal 't_a_79+slope' baseVal
+ t_a_80 baseVal 't_a_80+slope' peakVal
+ t_a_81 peakVal 't_a_81+slope' baseVal
+ t_a_82 baseVal 't_a_82+slope' peakVal
+ t_a_83 peakVal 't_a_83+slope' baseVal
+ t_a_84 baseVal 't_a_84+slope' peakVal
+ t_a_85 peakVal 't_a_85+slope' baseVal
+ t_a_86 baseVal 't_a_86+slope' peakVal
+ t_a_87 peakVal 't_a_87+slope' baseVal
+ t_a_88 baseVal 't_a_88+slope' peakVal
+ t_a_89 peakVal 't_a_89+slope' baseVal
+ t_a_90 baseVal 't_a_90+slope' peakVal
+ t_a_91 peakVal 't_a_91+slope' baseVal
+ t_a_92 baseVal 't_a_92+slope' peakVal
+ t_a_93 peakVal 't_a_93+slope' baseVal
+ t_a_94 baseVal 't_a_94+slope' peakVal
+ t_a_95 peakVal 't_a_95+slope' baseVal
+ t_a_96 baseVal 't_a_96+slope' peakVal
+ t_a_97 peakVal 't_a_97+slope' baseVal
+ t_a_98 baseVal 't_a_98+slope' peakVal
+ t_a_99 peakVal 't_a_99+slope' baseVal
+ t_a_100 baseVal 't_a_100+slope' peakVal
+ t_a_101 peakVal 't_a_101+slope' baseVal
+ t_a_102 baseVal 't_a_102+slope' peakVal
+ t_a_103 peakVal 't_a_103+slope' baseVal
+ t_a_104 baseVal 't_a_104+slope' peakVal
+ t_a_105 peakVal 't_a_105+slope' baseVal
+ t_a_106 baseVal 't_a_106+slope' peakVal
+ t_a_107 peakVal 't_a_107+slope' baseVal
+ t_a_108 baseVal 't_a_108+slope' peakVal
+ t_a_109 peakVal 't_a_109+slope' baseVal
+ t_a_110 baseVal 't_a_110+slope' peakVal
+ t_a_111 peakVal 't_a_111+slope' baseVal
+ t_a_112 baseVal 't_a_112+slope' peakVal
+ t_a_113 peakVal 't_a_113+slope' baseVal
+ t_a_114 baseVal 't_a_114+slope' peakVal
+ t_a_115 peakVal 't_a_115+slope' baseVal
+ t_a_116 baseVal 't_a_116+slope' peakVal
+ t_a_117 peakVal 't_a_117+slope' baseVal
+ t_a_118 baseVal 't_a_118+slope' peakVal
+ t_a_119 peakVal 't_a_119+slope' baseVal
+ t_a_120 baseVal 't_a_120+slope' peakVal
+ t_a_121 peakVal 't_a_121+slope' baseVal
+ t_a_122 baseVal 't_a_122+slope' peakVal
+ t_a_123 peakVal 't_a_123+slope' baseVal
+ t_a_124 baseVal 't_a_124+slope' peakVal
+ t_a_125 peakVal 't_a_125+slope' baseVal
+ t_a_126 baseVal 't_a_126+slope' peakVal
+ t_a_127 peakVal 't_a_127+slope' baseVal
+ t_a_128 baseVal 't_a_128+slope' peakVal
+ t_a_129 peakVal 't_a_129+slope' baseVal
+ t_a_130 baseVal 't_a_130+slope' peakVal
+ t_a_131 peakVal 't_a_131+slope' baseVal
+ t_a_132 baseVal 't_a_132+slope' peakVal
+ t_a_133 peakVal 't_a_133+slope' baseVal
+ t_a_134 baseVal 't_a_134+slope' peakVal
+ t_a_135 peakVal 't_a_135+slope' baseVal
+ t_a_136 baseVal 't_a_136+slope' peakVal
+ t_a_137 peakVal 't_a_137+slope' baseVal
+ t_a_138 baseVal 't_a_138+slope' peakVal
+ t_a_139 peakVal 't_a_139+slope' baseVal
+ t_a_140 baseVal 't_a_140+slope' peakVal
+ t_a_141 peakVal 't_a_141+slope' baseVal
+ t_a_142 baseVal 't_a_142+slope' peakVal
+ t_a_143 peakVal 't_a_143+slope' baseVal
+ t_a_144 baseVal 't_a_144+slope' peakVal
+ t_a_145 peakVal 't_a_145+slope' baseVal
+ t_a_146 baseVal 't_a_146+slope' peakVal
+ t_a_147 peakVal 't_a_147+slope' baseVal
+ t_a_148 baseVal 't_a_148+slope' peakVal
+ t_a_149 peakVal 't_a_149+slope' baseVal
+ t_a_150 baseVal 't_a_150+slope' peakVal
+ t_a_151 peakVal 't_a_151+slope' baseVal
+ t_a_152 baseVal 't_a_152+slope' peakVal
+ t_a_153 peakVal 't_a_153+slope' baseVal
+ t_a_154 baseVal 't_a_154+slope' peakVal
+ t_a_155 peakVal 't_a_155+slope' baseVal
+ t_a_156 baseVal 't_a_156+slope' peakVal
+ t_a_157 peakVal 't_a_157+slope' baseVal
+ t_a_158 baseVal 't_a_158+slope' peakVal
+ t_a_159 peakVal 't_a_159+slope' baseVal
+ t_a_160 baseVal 't_a_160+slope' peakVal
+ t_a_161 peakVal 't_a_161+slope' baseVal
+ t_a_162 baseVal 't_a_162+slope' peakVal
+ t_a_163 peakVal 't_a_163+slope' baseVal
+ t_a_164 baseVal 't_a_164+slope' peakVal
+ t_a_165 peakVal 't_a_165+slope' baseVal
+ t_a_166 baseVal 't_a_166+slope' peakVal
+ t_a_167 peakVal 't_a_167+slope' baseVal
+ t_a_168 baseVal 't_a_168+slope' peakVal
+ t_a_169 peakVal 't_a_169+slope' baseVal
+ t_a_170 baseVal 't_a_170+slope' peakVal
+ t_a_171 peakVal 't_a_171+slope' baseVal
+ t_a_172 baseVal 't_a_172+slope' peakVal
+ t_a_173 peakVal 't_a_173+slope' baseVal
+ t_a_174 baseVal 't_a_174+slope' peakVal
+ t_a_175 peakVal 't_a_175+slope' baseVal
+ t_a_176 baseVal 't_a_176+slope' peakVal
+ t_a_177 peakVal 't_a_177+slope' baseVal
+ t_a_178 baseVal 't_a_178+slope' peakVal
+ t_a_179 peakVal 't_a_179+slope' baseVal
+ t_a_180 baseVal 't_a_180+slope' peakVal
+ t_a_181 peakVal 't_a_181+slope' baseVal
+ t_a_182 baseVal 't_a_182+slope' peakVal
+ t_a_183 peakVal 't_a_183+slope' baseVal
+ t_a_184 baseVal 't_a_184+slope' peakVal
+ t_a_185 peakVal 't_a_185+slope' baseVal
+ t_a_186 baseVal 't_a_186+slope' peakVal
+ t_a_187 peakVal 't_a_187+slope' baseVal
+ t_a_188 baseVal 't_a_188+slope' peakVal
+ t_a_189 peakVal 't_a_189+slope' baseVal
+ t_a_190 baseVal 't_a_190+slope' peakVal
+ t_a_191 peakVal 't_a_191+slope' baseVal
+ t_a_192 baseVal 't_a_192+slope' peakVal
+ t_a_193 peakVal 't_a_193+slope' baseVal
+ t_a_194 baseVal 't_a_194+slope' peakVal
+ t_a_195 peakVal 't_a_195+slope' baseVal
+ t_a_196 baseVal 't_a_196+slope' peakVal
+ t_a_197 peakVal 't_a_197+slope' baseVal
+ t_a_198 baseVal 't_a_198+slope' peakVal
+ t_a_199 peakVal 't_a_199+slope' baseVal
+ t_a_200 baseVal 't_a_200+slope' peakVal
+ t_a_201 peakVal 't_a_201+slope' baseVal
+ t_a_202 baseVal 't_a_202+slope' peakVal
+ t_a_203 peakVal 't_a_203+slope' baseVal
+ t_a_204 baseVal 't_a_204+slope' peakVal
+ t_a_205 peakVal 't_a_205+slope' baseVal
+ t_a_206 baseVal 't_a_206+slope' peakVal
+ t_a_207 peakVal 't_a_207+slope' baseVal
+ t_a_208 baseVal 't_a_208+slope' peakVal
+ t_a_209 peakVal 't_a_209+slope' baseVal
+ t_a_210 baseVal 't_a_210+slope' peakVal
+ t_a_211 peakVal 't_a_211+slope' baseVal
+ t_a_212 baseVal 't_a_212+slope' peakVal
+ t_a_213 peakVal 't_a_213+slope' baseVal
+ t_a_214 baseVal 't_a_214+slope' peakVal
+ t_a_215 peakVal 't_a_215+slope' baseVal
+ t_a_216 baseVal 't_a_216+slope' peakVal
+ t_a_217 peakVal 't_a_217+slope' baseVal
+ t_a_218 baseVal 't_a_218+slope' peakVal
+ t_a_219 peakVal 't_a_219+slope' baseVal
+ t_a_220 baseVal 't_a_220+slope' peakVal
+ t_a_221 peakVal 't_a_221+slope' baseVal
+ t_a_222 baseVal 't_a_222+slope' peakVal
+ t_a_223 peakVal 't_a_223+slope' baseVal
+ t_a_224 baseVal 't_a_224+slope' peakVal
+ t_a_225 peakVal 't_a_225+slope' baseVal
+ t_a_226 baseVal 't_a_226+slope' peakVal
+ t_a_227 peakVal 't_a_227+slope' baseVal
+ t_a_228 baseVal 't_a_228+slope' peakVal
+ t_a_229 peakVal 't_a_229+slope' baseVal
+ t_a_230 baseVal 't_a_230+slope' peakVal
+ t_a_231 peakVal 't_a_231+slope' baseVal
+ t_a_232 baseVal 't_a_232+slope' peakVal
+ t_a_233 peakVal 't_a_233+slope' baseVal
+ t_a_234 baseVal 't_a_234+slope' peakVal
+ t_a_235 peakVal 't_a_235+slope' baseVal
+ t_a_236 baseVal 't_a_236+slope' peakVal
+ t_a_237 peakVal 't_a_237+slope' baseVal
+ t_a_238 baseVal 't_a_238+slope' peakVal
+ t_a_239 peakVal 't_a_239+slope' baseVal
+ t_a_240 baseVal 't_a_240+slope' peakVal
+ t_a_241 peakVal 't_a_241+slope' baseVal
+ t_a_242 baseVal 't_a_242+slope' peakVal
+ t_a_243 peakVal 't_a_243+slope' baseVal
+ t_a_244 baseVal 't_a_244+slope' peakVal
+ t_a_245 peakVal 't_a_245+slope' baseVal
+ t_a_246 baseVal 't_a_246+slope' peakVal
+ t_a_247 peakVal 't_a_247+slope' baseVal
+ t_a_248 baseVal 't_a_248+slope' peakVal
+ t_a_249 peakVal 't_a_249+slope' baseVal
+ t_a_250 baseVal 't_a_250+slope' peakVal
+ t_a_251 peakVal 't_a_251+slope' baseVal
+ t_a_252 baseVal 't_a_252+slope' peakVal
+ t_a_253 peakVal 't_a_253+slope' baseVal
+ t_a_254 baseVal 't_a_254+slope' peakVal
+ t_a_255 peakVal 't_a_255+slope' baseVal
+ t_a_256 baseVal 't_a_256+slope' peakVal
+ t_a_257 peakVal 't_a_257+slope' baseVal
+ t_a_258 baseVal 't_a_258+slope' peakVal
+ t_a_259 peakVal 't_a_259+slope' baseVal
+ t_a_260 baseVal 't_a_260+slope' peakVal
+ t_a_261 peakVal 't_a_261+slope' baseVal
+ t_a_262 baseVal 't_a_262+slope' peakVal
+ t_a_263 peakVal 't_a_263+slope' baseVal
+ t_a_264 baseVal 't_a_264+slope' peakVal
+ t_a_265 peakVal 't_a_265+slope' baseVal
+ t_a_266 baseVal 't_a_266+slope' peakVal
+ t_a_267 peakVal 't_a_267+slope' baseVal
+ t_a_268 baseVal 't_a_268+slope' peakVal
+ t_a_269 peakVal 't_a_269+slope' baseVal
+ t_a_270 baseVal 't_a_270+slope' peakVal
+ t_a_271 peakVal 't_a_271+slope' baseVal
+ t_a_272 baseVal 't_a_272+slope' peakVal
+ t_a_273 peakVal 't_a_273+slope' baseVal
+ t_a_274 baseVal 't_a_274+slope' peakVal
+ t_a_275 peakVal 't_a_275+slope' baseVal
+ t_a_276 baseVal 't_a_276+slope' peakVal
+ t_a_277 peakVal 't_a_277+slope' baseVal
+ t_a_278 baseVal 't_a_278+slope' peakVal
+ t_a_279 peakVal 't_a_279+slope' baseVal
+ t_a_280 baseVal 't_a_280+slope' peakVal
+ t_a_281 peakVal 't_a_281+slope' baseVal
+ t_a_282 baseVal 't_a_282+slope' peakVal
+ t_a_283 peakVal 't_a_283+slope' baseVal
+ t_a_284 baseVal 't_a_284+slope' peakVal
+ t_a_285 peakVal 't_a_285+slope' baseVal
+ t_a_286 baseVal 't_a_286+slope' peakVal
+ t_a_287 peakVal 't_a_287+slope' baseVal
+ t_a_288 baseVal 't_a_288+slope' peakVal
+ t_a_289 peakVal 't_a_289+slope' baseVal
+ t_a_290 baseVal 't_a_290+slope' peakVal
+ t_a_291 peakVal 't_a_291+slope' baseVal
+ t_a_292 baseVal 't_a_292+slope' peakVal
+ t_a_293 peakVal 't_a_293+slope' baseVal
+ t_a_294 baseVal 't_a_294+slope' peakVal
+ t_a_295 peakVal 't_a_295+slope' baseVal
+ t_a_296 baseVal 't_a_296+slope' peakVal
+ t_a_297 peakVal 't_a_297+slope' baseVal
+ t_a_298 baseVal 't_a_298+slope' peakVal
+ t_a_299 peakVal 't_a_299+slope' baseVal
+ t_a_300 baseVal 't_a_300+slope' peakVal
+ t_a_301 peakVal 't_a_301+slope' baseVal
+ t_a_302 baseVal 't_a_302+slope' peakVal
+ t_a_303 peakVal 't_a_303+slope' baseVal
+ t_a_304 baseVal 't_a_304+slope' peakVal
+ t_a_305 peakVal 't_a_305+slope' baseVal
+ t_a_306 baseVal 't_a_306+slope' peakVal
+ t_a_307 peakVal 't_a_307+slope' baseVal
+ t_a_308 baseVal 't_a_308+slope' peakVal
+ t_a_309 peakVal 't_a_309+slope' baseVal
+ t_a_310 baseVal 't_a_310+slope' peakVal
+ t_a_311 peakVal 't_a_311+slope' baseVal
+ t_a_312 baseVal 't_a_312+slope' peakVal
+ t_a_313 peakVal 't_a_313+slope' baseVal
+ t_a_314 baseVal 't_a_314+slope' peakVal
+ t_a_315 peakVal 't_a_315+slope' baseVal
+ t_a_316 baseVal 't_a_316+slope' peakVal
+ t_a_317 peakVal 't_a_317+slope' baseVal
+ t_a_318 baseVal 't_a_318+slope' peakVal
+ t_a_319 peakVal 't_a_319+slope' baseVal
+ t_a_320 baseVal 't_a_320+slope' peakVal
+ t_a_321 peakVal 't_a_321+slope' baseVal
+ t_a_322 baseVal 't_a_322+slope' peakVal
+ t_a_323 peakVal 't_a_323+slope' baseVal
+ t_a_324 baseVal 't_a_324+slope' peakVal
+ t_a_325 peakVal 't_a_325+slope' baseVal
+ t_a_326 baseVal 't_a_326+slope' peakVal
+ t_a_327 peakVal 't_a_327+slope' baseVal
+ t_a_328 baseVal 't_a_328+slope' peakVal
+ t_a_329 peakVal 't_a_329+slope' baseVal
+ t_a_330 baseVal 't_a_330+slope' peakVal
+ t_a_331 peakVal 't_a_331+slope' baseVal
+ t_a_332 baseVal 't_a_332+slope' peakVal
+ t_a_333 peakVal 't_a_333+slope' baseVal
+ t_a_334 baseVal 't_a_334+slope' peakVal
+ t_a_335 peakVal 't_a_335+slope' baseVal
+ t_a_336 baseVal 't_a_336+slope' peakVal
+ t_a_337 peakVal 't_a_337+slope' baseVal
+ t_a_338 baseVal 't_a_338+slope' peakVal
+ t_a_339 peakVal 't_a_339+slope' baseVal
+ t_a_340 baseVal 't_a_340+slope' peakVal
+ t_a_341 peakVal 't_a_341+slope' baseVal
+ t_a_342 baseVal 't_a_342+slope' peakVal
+ t_a_343 peakVal 't_a_343+slope' baseVal
+ t_a_344 baseVal 't_a_344+slope' peakVal
+ t_a_345 peakVal 't_a_345+slope' baseVal
+ t_a_346 baseVal 't_a_346+slope' peakVal
+ t_a_347 peakVal 't_a_347+slope' baseVal
+ t_a_348 baseVal 't_a_348+slope' peakVal
+ t_a_349 peakVal 't_a_349+slope' baseVal
+ t_a_350 baseVal 't_a_350+slope' peakVal
+ t_a_351 peakVal 't_a_351+slope' baseVal
+ t_a_352 baseVal 't_a_352+slope' peakVal
+ t_a_353 peakVal 't_a_353+slope' baseVal
+ t_a_354 baseVal 't_a_354+slope' peakVal
+ t_a_355 peakVal 't_a_355+slope' baseVal
+ t_a_356 baseVal 't_a_356+slope' peakVal
+ t_a_357 peakVal 't_a_357+slope' baseVal
+ t_a_358 baseVal 't_a_358+slope' peakVal
+ t_a_359 peakVal 't_a_359+slope' baseVal
+ t_a_360 baseVal 't_a_360+slope' peakVal
+ t_a_361 peakVal 't_a_361+slope' baseVal
+ t_a_362 baseVal 't_a_362+slope' peakVal
+ t_a_363 peakVal 't_a_363+slope' baseVal
+ t_a_364 baseVal 't_a_364+slope' peakVal
+ t_a_365 peakVal 't_a_365+slope' baseVal
+ t_a_366 baseVal 't_a_366+slope' peakVal
+ t_a_367 peakVal 't_a_367+slope' baseVal
+ t_a_368 baseVal 't_a_368+slope' peakVal
+ t_a_369 peakVal 't_a_369+slope' baseVal
+ t_a_370 baseVal 't_a_370+slope' peakVal
+ t_a_371 peakVal 't_a_371+slope' baseVal
+ t_a_372 baseVal 't_a_372+slope' peakVal
+ t_a_373 peakVal 't_a_373+slope' baseVal
+ t_a_374 baseVal 't_a_374+slope' peakVal
+ t_a_375 peakVal 't_a_375+slope' baseVal
+ t_a_376 baseVal 't_a_376+slope' peakVal
+ t_a_377 peakVal 't_a_377+slope' baseVal
+ t_a_378 baseVal 't_a_378+slope' peakVal
+ t_a_379 peakVal 't_a_379+slope' baseVal
+ t_a_380 baseVal 't_a_380+slope' peakVal
+ t_a_381 peakVal 't_a_381+slope' baseVal
+ t_a_382 baseVal 't_a_382+slope' peakVal
+ t_a_383 peakVal 't_a_383+slope' baseVal
+ t_a_384 baseVal 't_a_384+slope' peakVal
+ t_a_385 peakVal 't_a_385+slope' baseVal
+ t_a_386 baseVal 't_a_386+slope' peakVal
+ t_a_387 peakVal 't_a_387+slope' baseVal
+ t_a_388 baseVal 't_a_388+slope' peakVal
+ t_a_389 peakVal 't_a_389+slope' baseVal
+ t_a_390 baseVal 't_a_390+slope' peakVal
+ t_a_391 peakVal 't_a_391+slope' baseVal
+ t_a_392 baseVal 't_a_392+slope' peakVal
+ t_a_393 peakVal 't_a_393+slope' baseVal
+ t_a_394 baseVal 't_a_394+slope' peakVal
+ t_a_395 peakVal 't_a_395+slope' baseVal
+ t_a_396 baseVal 't_a_396+slope' peakVal
+ t_a_397 peakVal 't_a_397+slope' baseVal
+ t_a_398 baseVal 't_a_398+slope' peakVal
+ t_a_399 peakVal 't_a_399+slope' baseVal
+ t_a_400 baseVal 't_a_400+slope' peakVal
+ t_a_401 peakVal 't_a_401+slope' baseVal
+ t_a_402 baseVal 't_a_402+slope' peakVal
+ t_a_403 peakVal 't_a_403+slope' baseVal
+ t_a_404 baseVal 't_a_404+slope' peakVal
+ t_a_405 peakVal 't_a_405+slope' baseVal
+ t_a_406 baseVal 't_a_406+slope' peakVal
+ t_a_407 peakVal 't_a_407+slope' baseVal
+ t_a_408 baseVal 't_a_408+slope' peakVal
+ t_a_409 peakVal 't_a_409+slope' baseVal
+ t_a_410 baseVal 't_a_410+slope' peakVal
+ t_a_411 peakVal 't_a_411+slope' baseVal
+ t_a_412 baseVal 't_a_412+slope' peakVal
+ t_a_413 peakVal 't_a_413+slope' baseVal
+ t_a_414 baseVal 't_a_414+slope' peakVal
+ t_a_415 peakVal 't_a_415+slope' baseVal
+ t_a_416 baseVal 't_a_416+slope' peakVal
+ t_a_417 peakVal 't_a_417+slope' baseVal
+ t_a_418 baseVal 't_a_418+slope' peakVal
+ t_a_419 peakVal 't_a_419+slope' baseVal
+ t_a_420 baseVal 't_a_420+slope' peakVal
+ t_a_421 peakVal 't_a_421+slope' baseVal
+ t_a_422 baseVal 't_a_422+slope' peakVal
+ t_a_423 peakVal 't_a_423+slope' baseVal
+ t_a_424 baseVal 't_a_424+slope' peakVal
+ t_a_425 peakVal 't_a_425+slope' baseVal
+ t_a_426 baseVal 't_a_426+slope' peakVal
+ t_a_427 peakVal 't_a_427+slope' baseVal
+ t_a_428 baseVal 't_a_428+slope' peakVal
+ t_a_429 peakVal 't_a_429+slope' baseVal
+ t_a_430 baseVal 't_a_430+slope' peakVal
+ t_a_431 peakVal 't_a_431+slope' baseVal
+ t_a_432 baseVal 't_a_432+slope' peakVal
+ t_a_433 peakVal 't_a_433+slope' baseVal
+ t_a_434 baseVal 't_a_434+slope' peakVal
+ t_a_435 peakVal 't_a_435+slope' baseVal
+ t_a_436 baseVal 't_a_436+slope' peakVal
+ t_a_437 peakVal 't_a_437+slope' baseVal
+ t_a_438 baseVal 't_a_438+slope' peakVal
+ t_a_439 peakVal 't_a_439+slope' baseVal
+ t_a_440 baseVal 't_a_440+slope' peakVal
+ t_a_441 peakVal 't_a_441+slope' baseVal
+ t_a_442 baseVal 't_a_442+slope' peakVal
+ t_a_443 peakVal 't_a_443+slope' baseVal
+ t_a_444 baseVal 't_a_444+slope' peakVal
+ t_a_445 peakVal 't_a_445+slope' baseVal
+ t_a_446 baseVal 't_a_446+slope' peakVal
+ t_a_447 peakVal 't_a_447+slope' baseVal
+ t_a_448 baseVal 't_a_448+slope' peakVal
+ t_a_449 peakVal 't_a_449+slope' baseVal
+ t_a_450 baseVal 't_a_450+slope' peakVal
+ t_a_451 peakVal 't_a_451+slope' baseVal
+ t_a_452 baseVal 't_a_452+slope' peakVal
+ t_a_453 peakVal 't_a_453+slope' baseVal
+ t_a_454 baseVal 't_a_454+slope' peakVal
+ t_a_455 peakVal 't_a_455+slope' baseVal
+ t_a_456 baseVal 't_a_456+slope' peakVal
+ t_a_457 peakVal 't_a_457+slope' baseVal
+ t_a_458 baseVal 't_a_458+slope' peakVal
+ t_a_459 peakVal 't_a_459+slope' baseVal
+ t_a_460 baseVal 't_a_460+slope' peakVal
+ t_a_461 peakVal 't_a_461+slope' baseVal
+ t_a_462 baseVal 't_a_462+slope' peakVal
+ t_a_463 peakVal 't_a_463+slope' baseVal
+ t_a_464 baseVal 't_a_464+slope' peakVal
+ t_a_465 peakVal 't_a_465+slope' baseVal
+ t_a_466 baseVal 't_a_466+slope' peakVal
+ t_a_467 peakVal 't_a_467+slope' baseVal
+ t_a_468 baseVal 't_a_468+slope' peakVal
+ t_a_469 peakVal 't_a_469+slope' baseVal
+ t_a_470 baseVal 't_a_470+slope' peakVal
+ t_a_471 peakVal 't_a_471+slope' baseVal
+ t_a_472 baseVal 't_a_472+slope' peakVal
+ t_a_473 peakVal 't_a_473+slope' baseVal
+ t_a_474 baseVal 't_a_474+slope' peakVal
+ t_a_475 peakVal 't_a_475+slope' baseVal
+ t_a_476 baseVal 't_a_476+slope' peakVal
+ t_a_477 peakVal 't_a_477+slope' baseVal
+ t_a_478 baseVal 't_a_478+slope' peakVal
+ t_a_479 peakVal 't_a_479+slope' baseVal
+ t_a_480 baseVal 't_a_480+slope' peakVal
+ t_a_481 peakVal 't_a_481+slope' baseVal
+ t_a_482 baseVal 't_a_482+slope' peakVal
+ t_a_483 peakVal 't_a_483+slope' baseVal
+ t_a_484 baseVal 't_a_484+slope' peakVal
+ t_a_485 peakVal 't_a_485+slope' baseVal
+ t_a_486 baseVal 't_a_486+slope' peakVal
+ t_a_487 peakVal 't_a_487+slope' baseVal
+ t_a_488 baseVal 't_a_488+slope' peakVal
+ t_a_489 peakVal 't_a_489+slope' baseVal
+ t_a_490 baseVal 't_a_490+slope' peakVal
+ t_a_491 peakVal 't_a_491+slope' baseVal
+ t_a_492 baseVal 't_a_492+slope' peakVal
+ t_a_493 peakVal 't_a_493+slope' baseVal
+ t_a_494 baseVal 't_a_494+slope' peakVal
+ t_a_495 peakVal 't_a_495+slope' baseVal
+ t_a_496 baseVal 't_a_496+slope' peakVal
+ t_a_497 peakVal 't_a_497+slope' baseVal
+ t_a_498 baseVal 't_a_498+slope' peakVal
+ t_a_499 peakVal 't_a_499+slope' baseVal
+ t_a_500 baseVal 't_a_500+slope' peakVal
+ t_a_501 peakVal 't_a_501+slope' baseVal
+ t_a_502 baseVal 't_a_502+slope' peakVal
+ t_a_503 peakVal 't_a_503+slope' baseVal
+ t_a_504 baseVal 't_a_504+slope' peakVal
+ t_a_505 peakVal 't_a_505+slope' baseVal
+ t_a_506 baseVal 't_a_506+slope' peakVal
+ t_a_507 peakVal 't_a_507+slope' baseVal
+ t_a_508 baseVal 't_a_508+slope' peakVal
+ t_a_509 peakVal 't_a_509+slope' baseVal
+ t_a_510 baseVal 't_a_510+slope' peakVal
+ t_a_511 peakVal 't_a_511+slope' baseVal
+ t_a_512 baseVal 't_a_512+slope' peakVal
+ t_a_513 peakVal 't_a_513+slope' baseVal
+ t_a_514 baseVal 't_a_514+slope' peakVal
+ t_a_515 peakVal 't_a_515+slope' baseVal
+ t_a_516 baseVal 't_a_516+slope' peakVal
+ t_a_517 peakVal 't_a_517+slope' baseVal
+ t_a_518 baseVal 't_a_518+slope' peakVal
+ t_a_519 peakVal 't_a_519+slope' baseVal
+ t_a_520 baseVal 't_a_520+slope' peakVal
+ t_a_521 peakVal 't_a_521+slope' baseVal
+ t_a_522 baseVal 't_a_522+slope' peakVal
+ t_a_523 peakVal 't_a_523+slope' baseVal
+ t_a_524 baseVal 't_a_524+slope' peakVal
+ t_a_525 peakVal 't_a_525+slope' baseVal
+ t_a_526 baseVal 't_a_526+slope' peakVal
+ t_a_527 peakVal 't_a_527+slope' baseVal
+ t_a_528 baseVal 't_a_528+slope' peakVal
+ t_a_529 peakVal 't_a_529+slope' baseVal
+ t_a_530 baseVal 't_a_530+slope' peakVal
+ t_a_531 peakVal 't_a_531+slope' baseVal
+ t_a_532 baseVal 't_a_532+slope' peakVal
+ t_a_533 peakVal 't_a_533+slope' baseVal
+ t_a_534 baseVal 't_a_534+slope' peakVal
+ t_a_535 peakVal 't_a_535+slope' baseVal
+ t_a_536 baseVal 't_a_536+slope' peakVal
+ t_a_537 peakVal 't_a_537+slope' baseVal
+ t_a_538 baseVal 't_a_538+slope' peakVal
+ t_a_539 peakVal 't_a_539+slope' baseVal
+ t_a_540 baseVal 't_a_540+slope' peakVal
+ t_a_541 peakVal 't_a_541+slope' baseVal
+ t_a_542 baseVal 't_a_542+slope' peakVal
+ t_a_543 peakVal 't_a_543+slope' baseVal
+ t_a_544 baseVal 't_a_544+slope' peakVal
+ t_a_545 peakVal 't_a_545+slope' baseVal
+ t_a_546 baseVal 't_a_546+slope' peakVal
+ t_a_547 peakVal 't_a_547+slope' baseVal
+ t_a_548 baseVal 't_a_548+slope' peakVal
+ t_a_549 peakVal 't_a_549+slope' baseVal
+ t_a_550 baseVal 't_a_550+slope' peakVal
+ t_a_551 peakVal 't_a_551+slope' baseVal
+ t_a_552 baseVal 't_a_552+slope' peakVal
+ t_a_553 peakVal 't_a_553+slope' baseVal
+ t_a_554 baseVal 't_a_554+slope' peakVal
+ t_a_555 peakVal 't_a_555+slope' baseVal
+ t_a_556 baseVal 't_a_556+slope' peakVal
+ t_a_557 peakVal 't_a_557+slope' baseVal
+ t_a_558 baseVal 't_a_558+slope' peakVal
+ t_a_559 peakVal 't_a_559+slope' baseVal
+ t_a_560 baseVal 't_a_560+slope' peakVal
+ t_a_561 peakVal 't_a_561+slope' baseVal
+ t_a_562 baseVal 't_a_562+slope' peakVal
+ t_a_563 peakVal 't_a_563+slope' baseVal
+ t_a_564 baseVal 't_a_564+slope' peakVal
+ t_a_565 peakVal 't_a_565+slope' baseVal
+ t_a_566 baseVal 't_a_566+slope' peakVal
+ t_a_567 peakVal 't_a_567+slope' baseVal
+ t_a_568 baseVal 't_a_568+slope' peakVal
+ t_a_569 peakVal 't_a_569+slope' baseVal
+ t_a_570 baseVal 't_a_570+slope' peakVal
+ t_a_571 peakVal 't_a_571+slope' baseVal
+ t_a_572 baseVal 't_a_572+slope' peakVal
+ t_a_573 peakVal 't_a_573+slope' baseVal
+ t_a_574 baseVal 't_a_574+slope' peakVal
+ t_a_575 peakVal 't_a_575+slope' baseVal
+ t_a_576 baseVal 't_a_576+slope' peakVal
+ t_a_577 peakVal 't_a_577+slope' baseVal
+ t_a_578 baseVal 't_a_578+slope' peakVal
+ t_a_579 peakVal 't_a_579+slope' baseVal
+ t_a_580 baseVal 't_a_580+slope' peakVal
+ t_a_581 peakVal 't_a_581+slope' baseVal
+ t_a_582 baseVal 't_a_582+slope' peakVal
+ t_a_583 peakVal 't_a_583+slope' baseVal
+ t_a_584 baseVal 't_a_584+slope' peakVal
+ t_a_585 peakVal 't_a_585+slope' baseVal
+ t_a_586 baseVal 't_a_586+slope' peakVal
+ t_a_587 peakVal 't_a_587+slope' baseVal
+ t_a_588 baseVal 't_a_588+slope' peakVal
+ t_a_589 peakVal 't_a_589+slope' baseVal
+ t_a_590 baseVal 't_a_590+slope' peakVal
+ t_a_591 peakVal 't_a_591+slope' baseVal
+ t_a_592 baseVal 't_a_592+slope' peakVal
+ t_a_593 peakVal 't_a_593+slope' baseVal
+ t_a_594 baseVal 't_a_594+slope' peakVal
+ t_a_595 peakVal 't_a_595+slope' baseVal
+ t_a_596 baseVal 't_a_596+slope' peakVal
+ t_a_597 peakVal 't_a_597+slope' baseVal
+ t_a_598 baseVal 't_a_598+slope' peakVal
+ t_a_599 peakVal 't_a_599+slope' baseVal
+ t_a_600 baseVal 't_a_600+slope' peakVal
+ t_a_601 peakVal 't_a_601+slope' baseVal
+ t_a_602 baseVal 't_a_602+slope' peakVal
+ t_a_603 peakVal 't_a_603+slope' baseVal
+ t_a_604 baseVal 't_a_604+slope' peakVal
+ t_a_605 peakVal 't_a_605+slope' baseVal
+ t_a_606 baseVal 't_a_606+slope' peakVal
+ t_a_607 peakVal 't_a_607+slope' baseVal
+ t_a_608 baseVal 't_a_608+slope' peakVal
+ t_a_609 peakVal 't_a_609+slope' baseVal
+ t_a_610 baseVal 't_a_610+slope' peakVal
+ t_a_611 peakVal 't_a_611+slope' baseVal
+ t_a_612 baseVal 't_a_612+slope' peakVal
+ t_a_613 peakVal 't_a_613+slope' baseVal
+ t_a_614 baseVal 't_a_614+slope' peakVal
+ t_a_615 peakVal 't_a_615+slope' baseVal
+ t_a_616 baseVal 't_a_616+slope' peakVal
+ t_a_617 peakVal 't_a_617+slope' baseVal
+ t_a_618 baseVal 't_a_618+slope' peakVal
+ t_a_619 peakVal 't_a_619+slope' baseVal
+ t_a_620 baseVal 't_a_620+slope' peakVal
+ t_a_621 peakVal 't_a_621+slope' baseVal
+ t_a_622 baseVal 't_a_622+slope' peakVal
+ t_a_623 peakVal 't_a_623+slope' baseVal
+ t_a_624 baseVal 't_a_624+slope' peakVal
+ t_a_625 peakVal 't_a_625+slope' baseVal
+ t_a_626 baseVal 't_a_626+slope' peakVal
+ t_a_627 peakVal 't_a_627+slope' baseVal
+ t_a_628 baseVal 't_a_628+slope' peakVal
+ t_a_629 peakVal 't_a_629+slope' baseVal
+ t_a_630 baseVal 't_a_630+slope' peakVal
+ t_a_631 peakVal 't_a_631+slope' baseVal
+ t_a_632 baseVal 't_a_632+slope' peakVal
+ t_a_633 peakVal 't_a_633+slope' baseVal
+ t_a_634 baseVal 't_a_634+slope' peakVal
+ t_a_635 peakVal 't_a_635+slope' baseVal
+ t_a_636 baseVal 't_a_636+slope' peakVal
+ t_a_637 peakVal 't_a_637+slope' baseVal
+ t_a_638 baseVal 't_a_638+slope' peakVal
+ t_a_639 peakVal 't_a_639+slope' baseVal
+ t_a_640 baseVal 't_a_640+slope' peakVal
+ t_a_641 peakVal 't_a_641+slope' baseVal
+ t_a_642 baseVal 't_a_642+slope' peakVal
+ t_a_643 peakVal 't_a_643+slope' baseVal
+ t_a_644 baseVal 't_a_644+slope' peakVal
+ t_a_645 peakVal 't_a_645+slope' baseVal
+ t_a_646 baseVal 't_a_646+slope' peakVal
+ t_a_647 peakVal 't_a_647+slope' baseVal
+ t_a_648 baseVal 't_a_648+slope' peakVal
+ t_a_649 peakVal 't_a_649+slope' baseVal
+ t_a_650 baseVal 't_a_650+slope' peakVal
+ t_a_651 peakVal 't_a_651+slope' baseVal
+ t_a_652 baseVal 't_a_652+slope' peakVal
+ t_a_653 peakVal 't_a_653+slope' baseVal
+ t_a_654 baseVal 't_a_654+slope' peakVal
+ t_a_655 peakVal 't_a_655+slope' baseVal
+ t_a_656 baseVal 't_a_656+slope' peakVal
+ t_a_657 peakVal 't_a_657+slope' baseVal
+ t_a_658 baseVal 't_a_658+slope' peakVal
+ t_a_659 peakVal 't_a_659+slope' baseVal
+ t_a_660 baseVal 't_a_660+slope' peakVal
+ t_a_661 peakVal 't_a_661+slope' baseVal
+ t_a_662 baseVal 't_a_662+slope' peakVal
+ t_a_663 peakVal 't_a_663+slope' baseVal
+ t_a_664 baseVal 't_a_664+slope' peakVal
+ t_a_665 peakVal 't_a_665+slope' baseVal
+ t_a_666 baseVal 't_a_666+slope' peakVal
+ t_a_667 peakVal 't_a_667+slope' baseVal
+ t_a_668 baseVal 't_a_668+slope' peakVal
+ t_a_669 peakVal 't_a_669+slope' baseVal
+ t_a_670 baseVal 't_a_670+slope' peakVal
+ t_a_671 peakVal 't_a_671+slope' baseVal
+ t_a_672 baseVal 't_a_672+slope' peakVal
+ t_a_673 peakVal 't_a_673+slope' baseVal
+ t_a_674 baseVal 't_a_674+slope' peakVal
+ t_a_675 peakVal 't_a_675+slope' baseVal
+ t_a_676 baseVal 't_a_676+slope' peakVal
+ t_a_677 peakVal 't_a_677+slope' baseVal
+ t_a_678 baseVal 't_a_678+slope' peakVal
+ t_a_679 peakVal 't_a_679+slope' baseVal
+ t_a_680 baseVal 't_a_680+slope' peakVal
+ t_a_681 peakVal 't_a_681+slope' baseVal
+ t_a_682 baseVal 't_a_682+slope' peakVal
+ t_a_683 peakVal 't_a_683+slope' baseVal
+ t_a_684 baseVal 't_a_684+slope' peakVal
+ t_a_685 peakVal 't_a_685+slope' baseVal
+ t_a_686 baseVal 't_a_686+slope' peakVal
+ t_a_687 peakVal 't_a_687+slope' baseVal
+ t_a_688 baseVal 't_a_688+slope' peakVal
+ t_a_689 peakVal 't_a_689+slope' baseVal
+ t_a_690 baseVal 't_a_690+slope' peakVal
+ t_a_691 peakVal 't_a_691+slope' baseVal
+ t_a_692 baseVal 't_a_692+slope' peakVal
+ t_a_693 peakVal 't_a_693+slope' baseVal
+ t_a_694 baseVal 't_a_694+slope' peakVal
+ t_a_695 peakVal 't_a_695+slope' baseVal
+ t_a_696 baseVal 't_a_696+slope' peakVal
+ t_a_697 peakVal 't_a_697+slope' baseVal
+ t_a_698 baseVal 't_a_698+slope' peakVal
+ t_a_699 peakVal 't_a_699+slope' baseVal
+ t_a_700 baseVal 't_a_700+slope' peakVal
+ t_a_701 peakVal 't_a_701+slope' baseVal
+ t_a_702 baseVal 't_a_702+slope' peakVal
+ t_a_703 peakVal 't_a_703+slope' baseVal
+ t_a_704 baseVal 't_a_704+slope' peakVal
+ t_a_705 peakVal 't_a_705+slope' baseVal
+ t_a_706 baseVal 't_a_706+slope' peakVal
+ t_a_707 peakVal 't_a_707+slope' baseVal
+ t_a_708 baseVal 't_a_708+slope' peakVal
+ t_a_709 peakVal 't_a_709+slope' baseVal
+ t_a_710 baseVal 't_a_710+slope' peakVal
+ t_a_711 peakVal 't_a_711+slope' baseVal
+ t_a_712 baseVal 't_a_712+slope' peakVal
+ t_a_713 peakVal 't_a_713+slope' baseVal
+ t_a_714 baseVal 't_a_714+slope' peakVal
+ t_a_715 peakVal 't_a_715+slope' baseVal
+ t_a_716 baseVal 't_a_716+slope' peakVal
+ t_a_717 peakVal 't_a_717+slope' baseVal
+ t_a_718 baseVal 't_a_718+slope' peakVal
+ t_a_719 peakVal 't_a_719+slope' baseVal
+ t_a_720 baseVal 't_a_720+slope' peakVal
+ t_a_721 peakVal 't_a_721+slope' baseVal
+ t_a_722 baseVal 't_a_722+slope' peakVal
+ t_a_723 peakVal 't_a_723+slope' baseVal
+ t_a_724 baseVal 't_a_724+slope' peakVal
+ t_a_725 peakVal 't_a_725+slope' baseVal
+ t_a_726 baseVal 't_a_726+slope' peakVal
+ t_a_727 peakVal 't_a_727+slope' baseVal
+ t_a_728 baseVal 't_a_728+slope' peakVal
+ t_a_729 peakVal 't_a_729+slope' baseVal
+ t_a_730 baseVal 't_a_730+slope' peakVal
+ t_a_731 peakVal 't_a_731+slope' baseVal
+ t_a_732 baseVal 't_a_732+slope' peakVal
+ t_a_733 peakVal 't_a_733+slope' baseVal
+ t_a_734 baseVal 't_a_734+slope' peakVal
+ t_a_735 peakVal 't_a_735+slope' baseVal
+ t_a_736 baseVal 't_a_736+slope' peakVal
+ t_a_737 peakVal 't_a_737+slope' baseVal
+ t_a_738 baseVal 't_a_738+slope' peakVal
+ t_a_739 peakVal 't_a_739+slope' baseVal
+ t_a_740 baseVal 't_a_740+slope' peakVal
+ t_a_741 peakVal 't_a_741+slope' baseVal
+ t_a_742 baseVal 't_a_742+slope' peakVal
+ t_a_743 peakVal 't_a_743+slope' baseVal
+ t_a_744 baseVal 't_a_744+slope' peakVal
+ t_a_745 peakVal 't_a_745+slope' baseVal
+ t_a_746 baseVal 't_a_746+slope' peakVal
+ t_a_747 peakVal 't_a_747+slope' baseVal
+ t_a_748 baseVal 't_a_748+slope' peakVal
+ t_a_749 peakVal 't_a_749+slope' baseVal
+ t_a_750 baseVal 't_a_750+slope' peakVal
+ t_a_751 peakVal 't_a_751+slope' baseVal
+ t_a_752 baseVal 't_a_752+slope' peakVal
+ t_a_753 peakVal 't_a_753+slope' baseVal
+ t_a_754 baseVal 't_a_754+slope' peakVal
+ t_a_755 peakVal 't_a_755+slope' baseVal
+ t_a_756 baseVal 't_a_756+slope' peakVal
+ t_a_757 peakVal 't_a_757+slope' baseVal
+ t_a_758 baseVal 't_a_758+slope' peakVal
+ t_a_759 peakVal 't_a_759+slope' baseVal
+ t_a_760 baseVal 't_a_760+slope' peakVal
+ t_a_761 peakVal 't_a_761+slope' baseVal
+ t_a_762 baseVal 't_a_762+slope' peakVal
+ t_a_763 peakVal 't_a_763+slope' baseVal
+ t_a_764 baseVal 't_a_764+slope' peakVal
+ t_a_765 peakVal 't_a_765+slope' baseVal
+ t_a_766 baseVal 't_a_766+slope' peakVal
+ t_a_767 peakVal 't_a_767+slope' baseVal
+ t_a_768 baseVal 't_a_768+slope' peakVal
+ t_a_769 peakVal 't_a_769+slope' baseVal
+ t_a_770 baseVal 't_a_770+slope' peakVal
+ t_a_771 peakVal 't_a_771+slope' baseVal
+ t_a_772 baseVal 't_a_772+slope' peakVal
+ t_a_773 peakVal 't_a_773+slope' baseVal
+ t_a_774 baseVal 't_a_774+slope' peakVal
+ t_a_775 peakVal 't_a_775+slope' baseVal
+ t_a_776 baseVal 't_a_776+slope' peakVal
+ t_a_777 peakVal 't_a_777+slope' baseVal
+ t_a_778 baseVal 't_a_778+slope' peakVal
+ t_a_779 peakVal 't_a_779+slope' baseVal
+ t_a_780 baseVal 't_a_780+slope' peakVal
+ t_a_781 peakVal 't_a_781+slope' baseVal
+ t_a_782 baseVal 't_a_782+slope' peakVal
+ t_a_783 peakVal 't_a_783+slope' baseVal
+ t_a_784 baseVal 't_a_784+slope' peakVal
+ t_a_785 peakVal 't_a_785+slope' baseVal
+ t_a_786 baseVal 't_a_786+slope' peakVal
+ t_a_787 peakVal 't_a_787+slope' baseVal
+ t_a_788 baseVal 't_a_788+slope' peakVal
+ t_a_789 peakVal 't_a_789+slope' baseVal
+ t_a_790 baseVal 't_a_790+slope' peakVal
+ t_a_791 peakVal 't_a_791+slope' baseVal
+ t_a_792 baseVal 't_a_792+slope' peakVal
+ t_a_793 peakVal 't_a_793+slope' baseVal
+ t_a_794 baseVal 't_a_794+slope' peakVal
+ t_a_795 peakVal 't_a_795+slope' baseVal
+ t_a_796 baseVal 't_a_796+slope' peakVal
+ t_a_797 peakVal 't_a_797+slope' baseVal
+ t_a_798 baseVal 't_a_798+slope' peakVal
+ t_a_799 peakVal 't_a_799+slope' baseVal



VINB Input_B GND PWL 0ns baseVal t_init0 baseVal 't_init0+slope' peakVal t_init1 peakVal 't_init1+slope' baseVal
+ t_b_0 baseVal 't_b_0+slope' peakVal
+ t_b_1 peakVal 't_b_1+slope' baseVal
+ t_b_2 baseVal 't_b_2+slope' peakVal
+ t_b_3 peakVal 't_b_3+slope' baseVal
+ t_b_4 baseVal 't_b_4+slope' peakVal
+ t_b_5 peakVal 't_b_5+slope' baseVal
+ t_b_6 baseVal 't_b_6+slope' peakVal
+ t_b_7 peakVal 't_b_7+slope' baseVal
+ t_b_8 baseVal 't_b_8+slope' peakVal
+ t_b_9 peakVal 't_b_9+slope' baseVal
+ t_b_10 baseVal 't_b_10+slope' peakVal
+ t_b_11 peakVal 't_b_11+slope' baseVal
+ t_b_12 baseVal 't_b_12+slope' peakVal
+ t_b_13 peakVal 't_b_13+slope' baseVal
+ t_b_14 baseVal 't_b_14+slope' peakVal
+ t_b_15 peakVal 't_b_15+slope' baseVal
+ t_b_16 baseVal 't_b_16+slope' peakVal
+ t_b_17 peakVal 't_b_17+slope' baseVal
+ t_b_18 baseVal 't_b_18+slope' peakVal
+ t_b_19 peakVal 't_b_19+slope' baseVal
+ t_b_20 baseVal 't_b_20+slope' peakVal
+ t_b_21 peakVal 't_b_21+slope' baseVal
+ t_b_22 baseVal 't_b_22+slope' peakVal
+ t_b_23 peakVal 't_b_23+slope' baseVal
+ t_b_24 baseVal 't_b_24+slope' peakVal
+ t_b_25 peakVal 't_b_25+slope' baseVal
+ t_b_26 baseVal 't_b_26+slope' peakVal
+ t_b_27 peakVal 't_b_27+slope' baseVal
+ t_b_28 baseVal 't_b_28+slope' peakVal
+ t_b_29 peakVal 't_b_29+slope' baseVal
+ t_b_30 baseVal 't_b_30+slope' peakVal
+ t_b_31 peakVal 't_b_31+slope' baseVal
+ t_b_32 baseVal 't_b_32+slope' peakVal
+ t_b_33 peakVal 't_b_33+slope' baseVal
+ t_b_34 baseVal 't_b_34+slope' peakVal
+ t_b_35 peakVal 't_b_35+slope' baseVal
+ t_b_36 baseVal 't_b_36+slope' peakVal
+ t_b_37 peakVal 't_b_37+slope' baseVal
+ t_b_38 baseVal 't_b_38+slope' peakVal
+ t_b_39 peakVal 't_b_39+slope' baseVal
+ t_b_40 baseVal 't_b_40+slope' peakVal
+ t_b_41 peakVal 't_b_41+slope' baseVal
+ t_b_42 baseVal 't_b_42+slope' peakVal
+ t_b_43 peakVal 't_b_43+slope' baseVal
+ t_b_44 baseVal 't_b_44+slope' peakVal
+ t_b_45 peakVal 't_b_45+slope' baseVal
+ t_b_46 baseVal 't_b_46+slope' peakVal
+ t_b_47 peakVal 't_b_47+slope' baseVal
+ t_b_48 baseVal 't_b_48+slope' peakVal
+ t_b_49 peakVal 't_b_49+slope' baseVal
+ t_b_50 baseVal 't_b_50+slope' peakVal
+ t_b_51 peakVal 't_b_51+slope' baseVal
+ t_b_52 baseVal 't_b_52+slope' peakVal
+ t_b_53 peakVal 't_b_53+slope' baseVal
+ t_b_54 baseVal 't_b_54+slope' peakVal
+ t_b_55 peakVal 't_b_55+slope' baseVal
+ t_b_56 baseVal 't_b_56+slope' peakVal
+ t_b_57 peakVal 't_b_57+slope' baseVal
+ t_b_58 baseVal 't_b_58+slope' peakVal
+ t_b_59 peakVal 't_b_59+slope' baseVal
+ t_b_60 baseVal 't_b_60+slope' peakVal
+ t_b_61 peakVal 't_b_61+slope' baseVal
+ t_b_62 baseVal 't_b_62+slope' peakVal
+ t_b_63 peakVal 't_b_63+slope' baseVal
+ t_b_64 baseVal 't_b_64+slope' peakVal
+ t_b_65 peakVal 't_b_65+slope' baseVal
+ t_b_66 baseVal 't_b_66+slope' peakVal
+ t_b_67 peakVal 't_b_67+slope' baseVal
+ t_b_68 baseVal 't_b_68+slope' peakVal
+ t_b_69 peakVal 't_b_69+slope' baseVal
+ t_b_70 baseVal 't_b_70+slope' peakVal
+ t_b_71 peakVal 't_b_71+slope' baseVal
+ t_b_72 baseVal 't_b_72+slope' peakVal
+ t_b_73 peakVal 't_b_73+slope' baseVal
+ t_b_74 baseVal 't_b_74+slope' peakVal
+ t_b_75 peakVal 't_b_75+slope' baseVal
+ t_b_76 baseVal 't_b_76+slope' peakVal
+ t_b_77 peakVal 't_b_77+slope' baseVal
+ t_b_78 baseVal 't_b_78+slope' peakVal
+ t_b_79 peakVal 't_b_79+slope' baseVal
+ t_b_80 baseVal 't_b_80+slope' peakVal
+ t_b_81 peakVal 't_b_81+slope' baseVal
+ t_b_82 baseVal 't_b_82+slope' peakVal
+ t_b_83 peakVal 't_b_83+slope' baseVal
+ t_b_84 baseVal 't_b_84+slope' peakVal
+ t_b_85 peakVal 't_b_85+slope' baseVal
+ t_b_86 baseVal 't_b_86+slope' peakVal
+ t_b_87 peakVal 't_b_87+slope' baseVal
+ t_b_88 baseVal 't_b_88+slope' peakVal
+ t_b_89 peakVal 't_b_89+slope' baseVal
+ t_b_90 baseVal 't_b_90+slope' peakVal
+ t_b_91 peakVal 't_b_91+slope' baseVal
+ t_b_92 baseVal 't_b_92+slope' peakVal
+ t_b_93 peakVal 't_b_93+slope' baseVal
+ t_b_94 baseVal 't_b_94+slope' peakVal
+ t_b_95 peakVal 't_b_95+slope' baseVal
+ t_b_96 baseVal 't_b_96+slope' peakVal
+ t_b_97 peakVal 't_b_97+slope' baseVal
+ t_b_98 baseVal 't_b_98+slope' peakVal
+ t_b_99 peakVal 't_b_99+slope' baseVal
+ t_b_100 baseVal 't_b_100+slope' peakVal
+ t_b_101 peakVal 't_b_101+slope' baseVal
+ t_b_102 baseVal 't_b_102+slope' peakVal
+ t_b_103 peakVal 't_b_103+slope' baseVal
+ t_b_104 baseVal 't_b_104+slope' peakVal
+ t_b_105 peakVal 't_b_105+slope' baseVal
+ t_b_106 baseVal 't_b_106+slope' peakVal
+ t_b_107 peakVal 't_b_107+slope' baseVal
+ t_b_108 baseVal 't_b_108+slope' peakVal
+ t_b_109 peakVal 't_b_109+slope' baseVal
+ t_b_110 baseVal 't_b_110+slope' peakVal
+ t_b_111 peakVal 't_b_111+slope' baseVal
+ t_b_112 baseVal 't_b_112+slope' peakVal
+ t_b_113 peakVal 't_b_113+slope' baseVal
+ t_b_114 baseVal 't_b_114+slope' peakVal
+ t_b_115 peakVal 't_b_115+slope' baseVal
+ t_b_116 baseVal 't_b_116+slope' peakVal
+ t_b_117 peakVal 't_b_117+slope' baseVal
+ t_b_118 baseVal 't_b_118+slope' peakVal
+ t_b_119 peakVal 't_b_119+slope' baseVal
+ t_b_120 baseVal 't_b_120+slope' peakVal
+ t_b_121 peakVal 't_b_121+slope' baseVal
+ t_b_122 baseVal 't_b_122+slope' peakVal
+ t_b_123 peakVal 't_b_123+slope' baseVal
+ t_b_124 baseVal 't_b_124+slope' peakVal
+ t_b_125 peakVal 't_b_125+slope' baseVal
+ t_b_126 baseVal 't_b_126+slope' peakVal
+ t_b_127 peakVal 't_b_127+slope' baseVal
+ t_b_128 baseVal 't_b_128+slope' peakVal
+ t_b_129 peakVal 't_b_129+slope' baseVal
+ t_b_130 baseVal 't_b_130+slope' peakVal
+ t_b_131 peakVal 't_b_131+slope' baseVal
+ t_b_132 baseVal 't_b_132+slope' peakVal
+ t_b_133 peakVal 't_b_133+slope' baseVal
+ t_b_134 baseVal 't_b_134+slope' peakVal
+ t_b_135 peakVal 't_b_135+slope' baseVal
+ t_b_136 baseVal 't_b_136+slope' peakVal
+ t_b_137 peakVal 't_b_137+slope' baseVal
+ t_b_138 baseVal 't_b_138+slope' peakVal
+ t_b_139 peakVal 't_b_139+slope' baseVal
+ t_b_140 baseVal 't_b_140+slope' peakVal
+ t_b_141 peakVal 't_b_141+slope' baseVal
+ t_b_142 baseVal 't_b_142+slope' peakVal
+ t_b_143 peakVal 't_b_143+slope' baseVal
+ t_b_144 baseVal 't_b_144+slope' peakVal
+ t_b_145 peakVal 't_b_145+slope' baseVal
+ t_b_146 baseVal 't_b_146+slope' peakVal
+ t_b_147 peakVal 't_b_147+slope' baseVal
+ t_b_148 baseVal 't_b_148+slope' peakVal
+ t_b_149 peakVal 't_b_149+slope' baseVal
+ t_b_150 baseVal 't_b_150+slope' peakVal
+ t_b_151 peakVal 't_b_151+slope' baseVal
+ t_b_152 baseVal 't_b_152+slope' peakVal
+ t_b_153 peakVal 't_b_153+slope' baseVal
+ t_b_154 baseVal 't_b_154+slope' peakVal
+ t_b_155 peakVal 't_b_155+slope' baseVal
+ t_b_156 baseVal 't_b_156+slope' peakVal
+ t_b_157 peakVal 't_b_157+slope' baseVal
+ t_b_158 baseVal 't_b_158+slope' peakVal
+ t_b_159 peakVal 't_b_159+slope' baseVal
+ t_b_160 baseVal 't_b_160+slope' peakVal
+ t_b_161 peakVal 't_b_161+slope' baseVal
+ t_b_162 baseVal 't_b_162+slope' peakVal
+ t_b_163 peakVal 't_b_163+slope' baseVal
+ t_b_164 baseVal 't_b_164+slope' peakVal
+ t_b_165 peakVal 't_b_165+slope' baseVal
+ t_b_166 baseVal 't_b_166+slope' peakVal
+ t_b_167 peakVal 't_b_167+slope' baseVal
+ t_b_168 baseVal 't_b_168+slope' peakVal
+ t_b_169 peakVal 't_b_169+slope' baseVal
+ t_b_170 baseVal 't_b_170+slope' peakVal
+ t_b_171 peakVal 't_b_171+slope' baseVal
+ t_b_172 baseVal 't_b_172+slope' peakVal
+ t_b_173 peakVal 't_b_173+slope' baseVal
+ t_b_174 baseVal 't_b_174+slope' peakVal
+ t_b_175 peakVal 't_b_175+slope' baseVal
+ t_b_176 baseVal 't_b_176+slope' peakVal
+ t_b_177 peakVal 't_b_177+slope' baseVal
+ t_b_178 baseVal 't_b_178+slope' peakVal
+ t_b_179 peakVal 't_b_179+slope' baseVal
+ t_b_180 baseVal 't_b_180+slope' peakVal
+ t_b_181 peakVal 't_b_181+slope' baseVal
+ t_b_182 baseVal 't_b_182+slope' peakVal
+ t_b_183 peakVal 't_b_183+slope' baseVal
+ t_b_184 baseVal 't_b_184+slope' peakVal
+ t_b_185 peakVal 't_b_185+slope' baseVal
+ t_b_186 baseVal 't_b_186+slope' peakVal
+ t_b_187 peakVal 't_b_187+slope' baseVal
+ t_b_188 baseVal 't_b_188+slope' peakVal
+ t_b_189 peakVal 't_b_189+slope' baseVal
+ t_b_190 baseVal 't_b_190+slope' peakVal
+ t_b_191 peakVal 't_b_191+slope' baseVal
+ t_b_192 baseVal 't_b_192+slope' peakVal
+ t_b_193 peakVal 't_b_193+slope' baseVal
+ t_b_194 baseVal 't_b_194+slope' peakVal
+ t_b_195 peakVal 't_b_195+slope' baseVal
+ t_b_196 baseVal 't_b_196+slope' peakVal
+ t_b_197 peakVal 't_b_197+slope' baseVal
+ t_b_198 baseVal 't_b_198+slope' peakVal
+ t_b_199 peakVal 't_b_199+slope' baseVal
+ t_b_200 baseVal 't_b_200+slope' peakVal
+ t_b_201 peakVal 't_b_201+slope' baseVal
+ t_b_202 baseVal 't_b_202+slope' peakVal
+ t_b_203 peakVal 't_b_203+slope' baseVal
+ t_b_204 baseVal 't_b_204+slope' peakVal
+ t_b_205 peakVal 't_b_205+slope' baseVal
+ t_b_206 baseVal 't_b_206+slope' peakVal
+ t_b_207 peakVal 't_b_207+slope' baseVal
+ t_b_208 baseVal 't_b_208+slope' peakVal
+ t_b_209 peakVal 't_b_209+slope' baseVal
+ t_b_210 baseVal 't_b_210+slope' peakVal
+ t_b_211 peakVal 't_b_211+slope' baseVal
+ t_b_212 baseVal 't_b_212+slope' peakVal
+ t_b_213 peakVal 't_b_213+slope' baseVal
+ t_b_214 baseVal 't_b_214+slope' peakVal
+ t_b_215 peakVal 't_b_215+slope' baseVal
+ t_b_216 baseVal 't_b_216+slope' peakVal
+ t_b_217 peakVal 't_b_217+slope' baseVal
+ t_b_218 baseVal 't_b_218+slope' peakVal
+ t_b_219 peakVal 't_b_219+slope' baseVal
+ t_b_220 baseVal 't_b_220+slope' peakVal
+ t_b_221 peakVal 't_b_221+slope' baseVal
+ t_b_222 baseVal 't_b_222+slope' peakVal
+ t_b_223 peakVal 't_b_223+slope' baseVal
+ t_b_224 baseVal 't_b_224+slope' peakVal
+ t_b_225 peakVal 't_b_225+slope' baseVal
+ t_b_226 baseVal 't_b_226+slope' peakVal
+ t_b_227 peakVal 't_b_227+slope' baseVal
+ t_b_228 baseVal 't_b_228+slope' peakVal
+ t_b_229 peakVal 't_b_229+slope' baseVal
+ t_b_230 baseVal 't_b_230+slope' peakVal
+ t_b_231 peakVal 't_b_231+slope' baseVal
+ t_b_232 baseVal 't_b_232+slope' peakVal
+ t_b_233 peakVal 't_b_233+slope' baseVal
+ t_b_234 baseVal 't_b_234+slope' peakVal
+ t_b_235 peakVal 't_b_235+slope' baseVal
+ t_b_236 baseVal 't_b_236+slope' peakVal
+ t_b_237 peakVal 't_b_237+slope' baseVal
+ t_b_238 baseVal 't_b_238+slope' peakVal
+ t_b_239 peakVal 't_b_239+slope' baseVal
+ t_b_240 baseVal 't_b_240+slope' peakVal
+ t_b_241 peakVal 't_b_241+slope' baseVal
+ t_b_242 baseVal 't_b_242+slope' peakVal
+ t_b_243 peakVal 't_b_243+slope' baseVal
+ t_b_244 baseVal 't_b_244+slope' peakVal
+ t_b_245 peakVal 't_b_245+slope' baseVal
+ t_b_246 baseVal 't_b_246+slope' peakVal
+ t_b_247 peakVal 't_b_247+slope' baseVal
+ t_b_248 baseVal 't_b_248+slope' peakVal
+ t_b_249 peakVal 't_b_249+slope' baseVal
+ t_b_250 baseVal 't_b_250+slope' peakVal
+ t_b_251 peakVal 't_b_251+slope' baseVal
+ t_b_252 baseVal 't_b_252+slope' peakVal
+ t_b_253 peakVal 't_b_253+slope' baseVal
+ t_b_254 baseVal 't_b_254+slope' peakVal
+ t_b_255 peakVal 't_b_255+slope' baseVal
+ t_b_256 baseVal 't_b_256+slope' peakVal
+ t_b_257 peakVal 't_b_257+slope' baseVal
+ t_b_258 baseVal 't_b_258+slope' peakVal
+ t_b_259 peakVal 't_b_259+slope' baseVal
+ t_b_260 baseVal 't_b_260+slope' peakVal
+ t_b_261 peakVal 't_b_261+slope' baseVal
+ t_b_262 baseVal 't_b_262+slope' peakVal
+ t_b_263 peakVal 't_b_263+slope' baseVal
+ t_b_264 baseVal 't_b_264+slope' peakVal
+ t_b_265 peakVal 't_b_265+slope' baseVal
+ t_b_266 baseVal 't_b_266+slope' peakVal
+ t_b_267 peakVal 't_b_267+slope' baseVal
+ t_b_268 baseVal 't_b_268+slope' peakVal
+ t_b_269 peakVal 't_b_269+slope' baseVal
+ t_b_270 baseVal 't_b_270+slope' peakVal
+ t_b_271 peakVal 't_b_271+slope' baseVal
+ t_b_272 baseVal 't_b_272+slope' peakVal
+ t_b_273 peakVal 't_b_273+slope' baseVal
+ t_b_274 baseVal 't_b_274+slope' peakVal
+ t_b_275 peakVal 't_b_275+slope' baseVal
+ t_b_276 baseVal 't_b_276+slope' peakVal
+ t_b_277 peakVal 't_b_277+slope' baseVal
+ t_b_278 baseVal 't_b_278+slope' peakVal
+ t_b_279 peakVal 't_b_279+slope' baseVal
+ t_b_280 baseVal 't_b_280+slope' peakVal
+ t_b_281 peakVal 't_b_281+slope' baseVal
+ t_b_282 baseVal 't_b_282+slope' peakVal
+ t_b_283 peakVal 't_b_283+slope' baseVal
+ t_b_284 baseVal 't_b_284+slope' peakVal
+ t_b_285 peakVal 't_b_285+slope' baseVal
+ t_b_286 baseVal 't_b_286+slope' peakVal
+ t_b_287 peakVal 't_b_287+slope' baseVal
+ t_b_288 baseVal 't_b_288+slope' peakVal
+ t_b_289 peakVal 't_b_289+slope' baseVal
+ t_b_290 baseVal 't_b_290+slope' peakVal
+ t_b_291 peakVal 't_b_291+slope' baseVal
+ t_b_292 baseVal 't_b_292+slope' peakVal
+ t_b_293 peakVal 't_b_293+slope' baseVal
+ t_b_294 baseVal 't_b_294+slope' peakVal
+ t_b_295 peakVal 't_b_295+slope' baseVal
+ t_b_296 baseVal 't_b_296+slope' peakVal
+ t_b_297 peakVal 't_b_297+slope' baseVal
+ t_b_298 baseVal 't_b_298+slope' peakVal
+ t_b_299 peakVal 't_b_299+slope' baseVal
+ t_b_300 baseVal 't_b_300+slope' peakVal
+ t_b_301 peakVal 't_b_301+slope' baseVal
+ t_b_302 baseVal 't_b_302+slope' peakVal
+ t_b_303 peakVal 't_b_303+slope' baseVal
+ t_b_304 baseVal 't_b_304+slope' peakVal
+ t_b_305 peakVal 't_b_305+slope' baseVal
+ t_b_306 baseVal 't_b_306+slope' peakVal
+ t_b_307 peakVal 't_b_307+slope' baseVal
+ t_b_308 baseVal 't_b_308+slope' peakVal
+ t_b_309 peakVal 't_b_309+slope' baseVal
+ t_b_310 baseVal 't_b_310+slope' peakVal
+ t_b_311 peakVal 't_b_311+slope' baseVal
+ t_b_312 baseVal 't_b_312+slope' peakVal
+ t_b_313 peakVal 't_b_313+slope' baseVal
+ t_b_314 baseVal 't_b_314+slope' peakVal
+ t_b_315 peakVal 't_b_315+slope' baseVal
+ t_b_316 baseVal 't_b_316+slope' peakVal
+ t_b_317 peakVal 't_b_317+slope' baseVal
+ t_b_318 baseVal 't_b_318+slope' peakVal
+ t_b_319 peakVal 't_b_319+slope' baseVal
+ t_b_320 baseVal 't_b_320+slope' peakVal
+ t_b_321 peakVal 't_b_321+slope' baseVal
+ t_b_322 baseVal 't_b_322+slope' peakVal
+ t_b_323 peakVal 't_b_323+slope' baseVal
+ t_b_324 baseVal 't_b_324+slope' peakVal
+ t_b_325 peakVal 't_b_325+slope' baseVal
+ t_b_326 baseVal 't_b_326+slope' peakVal
+ t_b_327 peakVal 't_b_327+slope' baseVal
+ t_b_328 baseVal 't_b_328+slope' peakVal
+ t_b_329 peakVal 't_b_329+slope' baseVal
+ t_b_330 baseVal 't_b_330+slope' peakVal
+ t_b_331 peakVal 't_b_331+slope' baseVal
+ t_b_332 baseVal 't_b_332+slope' peakVal
+ t_b_333 peakVal 't_b_333+slope' baseVal
+ t_b_334 baseVal 't_b_334+slope' peakVal
+ t_b_335 peakVal 't_b_335+slope' baseVal
+ t_b_336 baseVal 't_b_336+slope' peakVal
+ t_b_337 peakVal 't_b_337+slope' baseVal
+ t_b_338 baseVal 't_b_338+slope' peakVal
+ t_b_339 peakVal 't_b_339+slope' baseVal
+ t_b_340 baseVal 't_b_340+slope' peakVal
+ t_b_341 peakVal 't_b_341+slope' baseVal
+ t_b_342 baseVal 't_b_342+slope' peakVal
+ t_b_343 peakVal 't_b_343+slope' baseVal
+ t_b_344 baseVal 't_b_344+slope' peakVal
+ t_b_345 peakVal 't_b_345+slope' baseVal
+ t_b_346 baseVal 't_b_346+slope' peakVal
+ t_b_347 peakVal 't_b_347+slope' baseVal
+ t_b_348 baseVal 't_b_348+slope' peakVal
+ t_b_349 peakVal 't_b_349+slope' baseVal
+ t_b_350 baseVal 't_b_350+slope' peakVal
+ t_b_351 peakVal 't_b_351+slope' baseVal
+ t_b_352 baseVal 't_b_352+slope' peakVal
+ t_b_353 peakVal 't_b_353+slope' baseVal
+ t_b_354 baseVal 't_b_354+slope' peakVal
+ t_b_355 peakVal 't_b_355+slope' baseVal
+ t_b_356 baseVal 't_b_356+slope' peakVal
+ t_b_357 peakVal 't_b_357+slope' baseVal
+ t_b_358 baseVal 't_b_358+slope' peakVal
+ t_b_359 peakVal 't_b_359+slope' baseVal
+ t_b_360 baseVal 't_b_360+slope' peakVal
+ t_b_361 peakVal 't_b_361+slope' baseVal
+ t_b_362 baseVal 't_b_362+slope' peakVal
+ t_b_363 peakVal 't_b_363+slope' baseVal
+ t_b_364 baseVal 't_b_364+slope' peakVal
+ t_b_365 peakVal 't_b_365+slope' baseVal
+ t_b_366 baseVal 't_b_366+slope' peakVal
+ t_b_367 peakVal 't_b_367+slope' baseVal
+ t_b_368 baseVal 't_b_368+slope' peakVal
+ t_b_369 peakVal 't_b_369+slope' baseVal
+ t_b_370 baseVal 't_b_370+slope' peakVal
+ t_b_371 peakVal 't_b_371+slope' baseVal
+ t_b_372 baseVal 't_b_372+slope' peakVal
+ t_b_373 peakVal 't_b_373+slope' baseVal
+ t_b_374 baseVal 't_b_374+slope' peakVal
+ t_b_375 peakVal 't_b_375+slope' baseVal
+ t_b_376 baseVal 't_b_376+slope' peakVal
+ t_b_377 peakVal 't_b_377+slope' baseVal
+ t_b_378 baseVal 't_b_378+slope' peakVal
+ t_b_379 peakVal 't_b_379+slope' baseVal
+ t_b_380 baseVal 't_b_380+slope' peakVal
+ t_b_381 peakVal 't_b_381+slope' baseVal
+ t_b_382 baseVal 't_b_382+slope' peakVal
+ t_b_383 peakVal 't_b_383+slope' baseVal
+ t_b_384 baseVal 't_b_384+slope' peakVal
+ t_b_385 peakVal 't_b_385+slope' baseVal
+ t_b_386 baseVal 't_b_386+slope' peakVal
+ t_b_387 peakVal 't_b_387+slope' baseVal
+ t_b_388 baseVal 't_b_388+slope' peakVal
+ t_b_389 peakVal 't_b_389+slope' baseVal
+ t_b_390 baseVal 't_b_390+slope' peakVal
+ t_b_391 peakVal 't_b_391+slope' baseVal
+ t_b_392 baseVal 't_b_392+slope' peakVal
+ t_b_393 peakVal 't_b_393+slope' baseVal
+ t_b_394 baseVal 't_b_394+slope' peakVal
+ t_b_395 peakVal 't_b_395+slope' baseVal
+ t_b_396 baseVal 't_b_396+slope' peakVal
+ t_b_397 peakVal 't_b_397+slope' baseVal
+ t_b_398 baseVal 't_b_398+slope' peakVal
+ t_b_399 peakVal 't_b_399+slope' baseVal
+ t_b_400 baseVal 't_b_400+slope' peakVal
+ t_b_401 peakVal 't_b_401+slope' baseVal
+ t_b_402 baseVal 't_b_402+slope' peakVal
+ t_b_403 peakVal 't_b_403+slope' baseVal
+ t_b_404 baseVal 't_b_404+slope' peakVal
+ t_b_405 peakVal 't_b_405+slope' baseVal
+ t_b_406 baseVal 't_b_406+slope' peakVal
+ t_b_407 peakVal 't_b_407+slope' baseVal
+ t_b_408 baseVal 't_b_408+slope' peakVal
+ t_b_409 peakVal 't_b_409+slope' baseVal
+ t_b_410 baseVal 't_b_410+slope' peakVal
+ t_b_411 peakVal 't_b_411+slope' baseVal
+ t_b_412 baseVal 't_b_412+slope' peakVal
+ t_b_413 peakVal 't_b_413+slope' baseVal
+ t_b_414 baseVal 't_b_414+slope' peakVal
+ t_b_415 peakVal 't_b_415+slope' baseVal
+ t_b_416 baseVal 't_b_416+slope' peakVal
+ t_b_417 peakVal 't_b_417+slope' baseVal
+ t_b_418 baseVal 't_b_418+slope' peakVal
+ t_b_419 peakVal 't_b_419+slope' baseVal
+ t_b_420 baseVal 't_b_420+slope' peakVal
+ t_b_421 peakVal 't_b_421+slope' baseVal
+ t_b_422 baseVal 't_b_422+slope' peakVal
+ t_b_423 peakVal 't_b_423+slope' baseVal
+ t_b_424 baseVal 't_b_424+slope' peakVal
+ t_b_425 peakVal 't_b_425+slope' baseVal
+ t_b_426 baseVal 't_b_426+slope' peakVal
+ t_b_427 peakVal 't_b_427+slope' baseVal
+ t_b_428 baseVal 't_b_428+slope' peakVal
+ t_b_429 peakVal 't_b_429+slope' baseVal
+ t_b_430 baseVal 't_b_430+slope' peakVal
+ t_b_431 peakVal 't_b_431+slope' baseVal
+ t_b_432 baseVal 't_b_432+slope' peakVal
+ t_b_433 peakVal 't_b_433+slope' baseVal
+ t_b_434 baseVal 't_b_434+slope' peakVal
+ t_b_435 peakVal 't_b_435+slope' baseVal
+ t_b_436 baseVal 't_b_436+slope' peakVal
+ t_b_437 peakVal 't_b_437+slope' baseVal
+ t_b_438 baseVal 't_b_438+slope' peakVal
+ t_b_439 peakVal 't_b_439+slope' baseVal
+ t_b_440 baseVal 't_b_440+slope' peakVal
+ t_b_441 peakVal 't_b_441+slope' baseVal
+ t_b_442 baseVal 't_b_442+slope' peakVal
+ t_b_443 peakVal 't_b_443+slope' baseVal
+ t_b_444 baseVal 't_b_444+slope' peakVal
+ t_b_445 peakVal 't_b_445+slope' baseVal
+ t_b_446 baseVal 't_b_446+slope' peakVal
+ t_b_447 peakVal 't_b_447+slope' baseVal
+ t_b_448 baseVal 't_b_448+slope' peakVal
+ t_b_449 peakVal 't_b_449+slope' baseVal
+ t_b_450 baseVal 't_b_450+slope' peakVal
+ t_b_451 peakVal 't_b_451+slope' baseVal
+ t_b_452 baseVal 't_b_452+slope' peakVal
+ t_b_453 peakVal 't_b_453+slope' baseVal
+ t_b_454 baseVal 't_b_454+slope' peakVal
+ t_b_455 peakVal 't_b_455+slope' baseVal
+ t_b_456 baseVal 't_b_456+slope' peakVal
+ t_b_457 peakVal 't_b_457+slope' baseVal
+ t_b_458 baseVal 't_b_458+slope' peakVal
+ t_b_459 peakVal 't_b_459+slope' baseVal
+ t_b_460 baseVal 't_b_460+slope' peakVal
+ t_b_461 peakVal 't_b_461+slope' baseVal
+ t_b_462 baseVal 't_b_462+slope' peakVal
+ t_b_463 peakVal 't_b_463+slope' baseVal
+ t_b_464 baseVal 't_b_464+slope' peakVal
+ t_b_465 peakVal 't_b_465+slope' baseVal
+ t_b_466 baseVal 't_b_466+slope' peakVal
+ t_b_467 peakVal 't_b_467+slope' baseVal
+ t_b_468 baseVal 't_b_468+slope' peakVal
+ t_b_469 peakVal 't_b_469+slope' baseVal
+ t_b_470 baseVal 't_b_470+slope' peakVal
+ t_b_471 peakVal 't_b_471+slope' baseVal
+ t_b_472 baseVal 't_b_472+slope' peakVal
+ t_b_473 peakVal 't_b_473+slope' baseVal
+ t_b_474 baseVal 't_b_474+slope' peakVal
+ t_b_475 peakVal 't_b_475+slope' baseVal
+ t_b_476 baseVal 't_b_476+slope' peakVal
+ t_b_477 peakVal 't_b_477+slope' baseVal
+ t_b_478 baseVal 't_b_478+slope' peakVal
+ t_b_479 peakVal 't_b_479+slope' baseVal
+ t_b_480 baseVal 't_b_480+slope' peakVal
+ t_b_481 peakVal 't_b_481+slope' baseVal
+ t_b_482 baseVal 't_b_482+slope' peakVal
+ t_b_483 peakVal 't_b_483+slope' baseVal
+ t_b_484 baseVal 't_b_484+slope' peakVal
+ t_b_485 peakVal 't_b_485+slope' baseVal
+ t_b_486 baseVal 't_b_486+slope' peakVal
+ t_b_487 peakVal 't_b_487+slope' baseVal
+ t_b_488 baseVal 't_b_488+slope' peakVal
+ t_b_489 peakVal 't_b_489+slope' baseVal
+ t_b_490 baseVal 't_b_490+slope' peakVal
+ t_b_491 peakVal 't_b_491+slope' baseVal
+ t_b_492 baseVal 't_b_492+slope' peakVal
+ t_b_493 peakVal 't_b_493+slope' baseVal
+ t_b_494 baseVal 't_b_494+slope' peakVal
+ t_b_495 peakVal 't_b_495+slope' baseVal
+ t_b_496 baseVal 't_b_496+slope' peakVal
+ t_b_497 peakVal 't_b_497+slope' baseVal
+ t_b_498 baseVal 't_b_498+slope' peakVal
+ t_b_499 peakVal 't_b_499+slope' baseVal
+ t_b_500 baseVal 't_b_500+slope' peakVal
+ t_b_501 peakVal 't_b_501+slope' baseVal
+ t_b_502 baseVal 't_b_502+slope' peakVal
+ t_b_503 peakVal 't_b_503+slope' baseVal
+ t_b_504 baseVal 't_b_504+slope' peakVal
+ t_b_505 peakVal 't_b_505+slope' baseVal
+ t_b_506 baseVal 't_b_506+slope' peakVal
+ t_b_507 peakVal 't_b_507+slope' baseVal
+ t_b_508 baseVal 't_b_508+slope' peakVal
+ t_b_509 peakVal 't_b_509+slope' baseVal
+ t_b_510 baseVal 't_b_510+slope' peakVal
+ t_b_511 peakVal 't_b_511+slope' baseVal
+ t_b_512 baseVal 't_b_512+slope' peakVal
+ t_b_513 peakVal 't_b_513+slope' baseVal
+ t_b_514 baseVal 't_b_514+slope' peakVal
+ t_b_515 peakVal 't_b_515+slope' baseVal
+ t_b_516 baseVal 't_b_516+slope' peakVal
+ t_b_517 peakVal 't_b_517+slope' baseVal
+ t_b_518 baseVal 't_b_518+slope' peakVal
+ t_b_519 peakVal 't_b_519+slope' baseVal
+ t_b_520 baseVal 't_b_520+slope' peakVal
+ t_b_521 peakVal 't_b_521+slope' baseVal
+ t_b_522 baseVal 't_b_522+slope' peakVal
+ t_b_523 peakVal 't_b_523+slope' baseVal
+ t_b_524 baseVal 't_b_524+slope' peakVal
+ t_b_525 peakVal 't_b_525+slope' baseVal
+ t_b_526 baseVal 't_b_526+slope' peakVal
+ t_b_527 peakVal 't_b_527+slope' baseVal
+ t_b_528 baseVal 't_b_528+slope' peakVal
+ t_b_529 peakVal 't_b_529+slope' baseVal
+ t_b_530 baseVal 't_b_530+slope' peakVal
+ t_b_531 peakVal 't_b_531+slope' baseVal
+ t_b_532 baseVal 't_b_532+slope' peakVal
+ t_b_533 peakVal 't_b_533+slope' baseVal
+ t_b_534 baseVal 't_b_534+slope' peakVal
+ t_b_535 peakVal 't_b_535+slope' baseVal
+ t_b_536 baseVal 't_b_536+slope' peakVal
+ t_b_537 peakVal 't_b_537+slope' baseVal
+ t_b_538 baseVal 't_b_538+slope' peakVal
+ t_b_539 peakVal 't_b_539+slope' baseVal
+ t_b_540 baseVal 't_b_540+slope' peakVal
+ t_b_541 peakVal 't_b_541+slope' baseVal
+ t_b_542 baseVal 't_b_542+slope' peakVal
+ t_b_543 peakVal 't_b_543+slope' baseVal
+ t_b_544 baseVal 't_b_544+slope' peakVal
+ t_b_545 peakVal 't_b_545+slope' baseVal
+ t_b_546 baseVal 't_b_546+slope' peakVal
+ t_b_547 peakVal 't_b_547+slope' baseVal
+ t_b_548 baseVal 't_b_548+slope' peakVal
+ t_b_549 peakVal 't_b_549+slope' baseVal
+ t_b_550 baseVal 't_b_550+slope' peakVal
+ t_b_551 peakVal 't_b_551+slope' baseVal
+ t_b_552 baseVal 't_b_552+slope' peakVal
+ t_b_553 peakVal 't_b_553+slope' baseVal
+ t_b_554 baseVal 't_b_554+slope' peakVal
+ t_b_555 peakVal 't_b_555+slope' baseVal
+ t_b_556 baseVal 't_b_556+slope' peakVal
+ t_b_557 peakVal 't_b_557+slope' baseVal
+ t_b_558 baseVal 't_b_558+slope' peakVal
+ t_b_559 peakVal 't_b_559+slope' baseVal
+ t_b_560 baseVal 't_b_560+slope' peakVal
+ t_b_561 peakVal 't_b_561+slope' baseVal
+ t_b_562 baseVal 't_b_562+slope' peakVal
+ t_b_563 peakVal 't_b_563+slope' baseVal
+ t_b_564 baseVal 't_b_564+slope' peakVal
+ t_b_565 peakVal 't_b_565+slope' baseVal
+ t_b_566 baseVal 't_b_566+slope' peakVal
+ t_b_567 peakVal 't_b_567+slope' baseVal
+ t_b_568 baseVal 't_b_568+slope' peakVal
+ t_b_569 peakVal 't_b_569+slope' baseVal
+ t_b_570 baseVal 't_b_570+slope' peakVal
+ t_b_571 peakVal 't_b_571+slope' baseVal
+ t_b_572 baseVal 't_b_572+slope' peakVal
+ t_b_573 peakVal 't_b_573+slope' baseVal
+ t_b_574 baseVal 't_b_574+slope' peakVal
+ t_b_575 peakVal 't_b_575+slope' baseVal
+ t_b_576 baseVal 't_b_576+slope' peakVal
+ t_b_577 peakVal 't_b_577+slope' baseVal
+ t_b_578 baseVal 't_b_578+slope' peakVal
+ t_b_579 peakVal 't_b_579+slope' baseVal
+ t_b_580 baseVal 't_b_580+slope' peakVal
+ t_b_581 peakVal 't_b_581+slope' baseVal
+ t_b_582 baseVal 't_b_582+slope' peakVal
+ t_b_583 peakVal 't_b_583+slope' baseVal
+ t_b_584 baseVal 't_b_584+slope' peakVal
+ t_b_585 peakVal 't_b_585+slope' baseVal
+ t_b_586 baseVal 't_b_586+slope' peakVal
+ t_b_587 peakVal 't_b_587+slope' baseVal
+ t_b_588 baseVal 't_b_588+slope' peakVal
+ t_b_589 peakVal 't_b_589+slope' baseVal
+ t_b_590 baseVal 't_b_590+slope' peakVal
+ t_b_591 peakVal 't_b_591+slope' baseVal
+ t_b_592 baseVal 't_b_592+slope' peakVal
+ t_b_593 peakVal 't_b_593+slope' baseVal
+ t_b_594 baseVal 't_b_594+slope' peakVal
+ t_b_595 peakVal 't_b_595+slope' baseVal
+ t_b_596 baseVal 't_b_596+slope' peakVal
+ t_b_597 peakVal 't_b_597+slope' baseVal
+ t_b_598 baseVal 't_b_598+slope' peakVal
+ t_b_599 peakVal 't_b_599+slope' baseVal
+ t_b_600 baseVal 't_b_600+slope' peakVal
+ t_b_601 peakVal 't_b_601+slope' baseVal
+ t_b_602 baseVal 't_b_602+slope' peakVal
+ t_b_603 peakVal 't_b_603+slope' baseVal
+ t_b_604 baseVal 't_b_604+slope' peakVal
+ t_b_605 peakVal 't_b_605+slope' baseVal
+ t_b_606 baseVal 't_b_606+slope' peakVal
+ t_b_607 peakVal 't_b_607+slope' baseVal
+ t_b_608 baseVal 't_b_608+slope' peakVal
+ t_b_609 peakVal 't_b_609+slope' baseVal
+ t_b_610 baseVal 't_b_610+slope' peakVal
+ t_b_611 peakVal 't_b_611+slope' baseVal
+ t_b_612 baseVal 't_b_612+slope' peakVal
+ t_b_613 peakVal 't_b_613+slope' baseVal
+ t_b_614 baseVal 't_b_614+slope' peakVal
+ t_b_615 peakVal 't_b_615+slope' baseVal
+ t_b_616 baseVal 't_b_616+slope' peakVal
+ t_b_617 peakVal 't_b_617+slope' baseVal
+ t_b_618 baseVal 't_b_618+slope' peakVal
+ t_b_619 peakVal 't_b_619+slope' baseVal
+ t_b_620 baseVal 't_b_620+slope' peakVal
+ t_b_621 peakVal 't_b_621+slope' baseVal
+ t_b_622 baseVal 't_b_622+slope' peakVal
+ t_b_623 peakVal 't_b_623+slope' baseVal
+ t_b_624 baseVal 't_b_624+slope' peakVal
+ t_b_625 peakVal 't_b_625+slope' baseVal
+ t_b_626 baseVal 't_b_626+slope' peakVal
+ t_b_627 peakVal 't_b_627+slope' baseVal
+ t_b_628 baseVal 't_b_628+slope' peakVal
+ t_b_629 peakVal 't_b_629+slope' baseVal
+ t_b_630 baseVal 't_b_630+slope' peakVal
+ t_b_631 peakVal 't_b_631+slope' baseVal
+ t_b_632 baseVal 't_b_632+slope' peakVal
+ t_b_633 peakVal 't_b_633+slope' baseVal
+ t_b_634 baseVal 't_b_634+slope' peakVal
+ t_b_635 peakVal 't_b_635+slope' baseVal
+ t_b_636 baseVal 't_b_636+slope' peakVal
+ t_b_637 peakVal 't_b_637+slope' baseVal
+ t_b_638 baseVal 't_b_638+slope' peakVal
+ t_b_639 peakVal 't_b_639+slope' baseVal
+ t_b_640 baseVal 't_b_640+slope' peakVal
+ t_b_641 peakVal 't_b_641+slope' baseVal
+ t_b_642 baseVal 't_b_642+slope' peakVal
+ t_b_643 peakVal 't_b_643+slope' baseVal
+ t_b_644 baseVal 't_b_644+slope' peakVal
+ t_b_645 peakVal 't_b_645+slope' baseVal
+ t_b_646 baseVal 't_b_646+slope' peakVal
+ t_b_647 peakVal 't_b_647+slope' baseVal
+ t_b_648 baseVal 't_b_648+slope' peakVal
+ t_b_649 peakVal 't_b_649+slope' baseVal
+ t_b_650 baseVal 't_b_650+slope' peakVal
+ t_b_651 peakVal 't_b_651+slope' baseVal
+ t_b_652 baseVal 't_b_652+slope' peakVal
+ t_b_653 peakVal 't_b_653+slope' baseVal
+ t_b_654 baseVal 't_b_654+slope' peakVal
+ t_b_655 peakVal 't_b_655+slope' baseVal
+ t_b_656 baseVal 't_b_656+slope' peakVal
+ t_b_657 peakVal 't_b_657+slope' baseVal
+ t_b_658 baseVal 't_b_658+slope' peakVal
+ t_b_659 peakVal 't_b_659+slope' baseVal
+ t_b_660 baseVal 't_b_660+slope' peakVal
+ t_b_661 peakVal 't_b_661+slope' baseVal
+ t_b_662 baseVal 't_b_662+slope' peakVal
+ t_b_663 peakVal 't_b_663+slope' baseVal
+ t_b_664 baseVal 't_b_664+slope' peakVal
+ t_b_665 peakVal 't_b_665+slope' baseVal
+ t_b_666 baseVal 't_b_666+slope' peakVal
+ t_b_667 peakVal 't_b_667+slope' baseVal
+ t_b_668 baseVal 't_b_668+slope' peakVal
+ t_b_669 peakVal 't_b_669+slope' baseVal
+ t_b_670 baseVal 't_b_670+slope' peakVal
+ t_b_671 peakVal 't_b_671+slope' baseVal
+ t_b_672 baseVal 't_b_672+slope' peakVal
+ t_b_673 peakVal 't_b_673+slope' baseVal
+ t_b_674 baseVal 't_b_674+slope' peakVal
+ t_b_675 peakVal 't_b_675+slope' baseVal
+ t_b_676 baseVal 't_b_676+slope' peakVal
+ t_b_677 peakVal 't_b_677+slope' baseVal
+ t_b_678 baseVal 't_b_678+slope' peakVal
+ t_b_679 peakVal 't_b_679+slope' baseVal
+ t_b_680 baseVal 't_b_680+slope' peakVal
+ t_b_681 peakVal 't_b_681+slope' baseVal
+ t_b_682 baseVal 't_b_682+slope' peakVal
+ t_b_683 peakVal 't_b_683+slope' baseVal
+ t_b_684 baseVal 't_b_684+slope' peakVal
+ t_b_685 peakVal 't_b_685+slope' baseVal
+ t_b_686 baseVal 't_b_686+slope' peakVal
+ t_b_687 peakVal 't_b_687+slope' baseVal
+ t_b_688 baseVal 't_b_688+slope' peakVal
+ t_b_689 peakVal 't_b_689+slope' baseVal
+ t_b_690 baseVal 't_b_690+slope' peakVal
+ t_b_691 peakVal 't_b_691+slope' baseVal
+ t_b_692 baseVal 't_b_692+slope' peakVal
+ t_b_693 peakVal 't_b_693+slope' baseVal
+ t_b_694 baseVal 't_b_694+slope' peakVal
+ t_b_695 peakVal 't_b_695+slope' baseVal
+ t_b_696 baseVal 't_b_696+slope' peakVal
+ t_b_697 peakVal 't_b_697+slope' baseVal
+ t_b_698 baseVal 't_b_698+slope' peakVal
+ t_b_699 peakVal 't_b_699+slope' baseVal
+ t_b_700 baseVal 't_b_700+slope' peakVal
+ t_b_701 peakVal 't_b_701+slope' baseVal
+ t_b_702 baseVal 't_b_702+slope' peakVal
+ t_b_703 peakVal 't_b_703+slope' baseVal
+ t_b_704 baseVal 't_b_704+slope' peakVal
+ t_b_705 peakVal 't_b_705+slope' baseVal
+ t_b_706 baseVal 't_b_706+slope' peakVal
+ t_b_707 peakVal 't_b_707+slope' baseVal
+ t_b_708 baseVal 't_b_708+slope' peakVal
+ t_b_709 peakVal 't_b_709+slope' baseVal
+ t_b_710 baseVal 't_b_710+slope' peakVal
+ t_b_711 peakVal 't_b_711+slope' baseVal
+ t_b_712 baseVal 't_b_712+slope' peakVal
+ t_b_713 peakVal 't_b_713+slope' baseVal
+ t_b_714 baseVal 't_b_714+slope' peakVal
+ t_b_715 peakVal 't_b_715+slope' baseVal
+ t_b_716 baseVal 't_b_716+slope' peakVal
+ t_b_717 peakVal 't_b_717+slope' baseVal
+ t_b_718 baseVal 't_b_718+slope' peakVal
+ t_b_719 peakVal 't_b_719+slope' baseVal
+ t_b_720 baseVal 't_b_720+slope' peakVal
+ t_b_721 peakVal 't_b_721+slope' baseVal
+ t_b_722 baseVal 't_b_722+slope' peakVal
+ t_b_723 peakVal 't_b_723+slope' baseVal
+ t_b_724 baseVal 't_b_724+slope' peakVal
+ t_b_725 peakVal 't_b_725+slope' baseVal
+ t_b_726 baseVal 't_b_726+slope' peakVal
+ t_b_727 peakVal 't_b_727+slope' baseVal
+ t_b_728 baseVal 't_b_728+slope' peakVal
+ t_b_729 peakVal 't_b_729+slope' baseVal
+ t_b_730 baseVal 't_b_730+slope' peakVal
+ t_b_731 peakVal 't_b_731+slope' baseVal
+ t_b_732 baseVal 't_b_732+slope' peakVal
+ t_b_733 peakVal 't_b_733+slope' baseVal
+ t_b_734 baseVal 't_b_734+slope' peakVal
+ t_b_735 peakVal 't_b_735+slope' baseVal
+ t_b_736 baseVal 't_b_736+slope' peakVal
+ t_b_737 peakVal 't_b_737+slope' baseVal
+ t_b_738 baseVal 't_b_738+slope' peakVal
+ t_b_739 peakVal 't_b_739+slope' baseVal
+ t_b_740 baseVal 't_b_740+slope' peakVal
+ t_b_741 peakVal 't_b_741+slope' baseVal
+ t_b_742 baseVal 't_b_742+slope' peakVal
+ t_b_743 peakVal 't_b_743+slope' baseVal
+ t_b_744 baseVal 't_b_744+slope' peakVal
+ t_b_745 peakVal 't_b_745+slope' baseVal
+ t_b_746 baseVal 't_b_746+slope' peakVal
+ t_b_747 peakVal 't_b_747+slope' baseVal
+ t_b_748 baseVal 't_b_748+slope' peakVal
+ t_b_749 peakVal 't_b_749+slope' baseVal
+ t_b_750 baseVal 't_b_750+slope' peakVal
+ t_b_751 peakVal 't_b_751+slope' baseVal
+ t_b_752 baseVal 't_b_752+slope' peakVal
+ t_b_753 peakVal 't_b_753+slope' baseVal
+ t_b_754 baseVal 't_b_754+slope' peakVal
+ t_b_755 peakVal 't_b_755+slope' baseVal
+ t_b_756 baseVal 't_b_756+slope' peakVal
+ t_b_757 peakVal 't_b_757+slope' baseVal
+ t_b_758 baseVal 't_b_758+slope' peakVal
+ t_b_759 peakVal 't_b_759+slope' baseVal
+ t_b_760 baseVal 't_b_760+slope' peakVal
+ t_b_761 peakVal 't_b_761+slope' baseVal
+ t_b_762 baseVal 't_b_762+slope' peakVal
+ t_b_763 peakVal 't_b_763+slope' baseVal
+ t_b_764 baseVal 't_b_764+slope' peakVal
+ t_b_765 peakVal 't_b_765+slope' baseVal
+ t_b_766 baseVal 't_b_766+slope' peakVal
+ t_b_767 peakVal 't_b_767+slope' baseVal
+ t_b_768 baseVal 't_b_768+slope' peakVal
+ t_b_769 peakVal 't_b_769+slope' baseVal
+ t_b_770 baseVal 't_b_770+slope' peakVal
+ t_b_771 peakVal 't_b_771+slope' baseVal
+ t_b_772 baseVal 't_b_772+slope' peakVal
+ t_b_773 peakVal 't_b_773+slope' baseVal
+ t_b_774 baseVal 't_b_774+slope' peakVal
+ t_b_775 peakVal 't_b_775+slope' baseVal
+ t_b_776 baseVal 't_b_776+slope' peakVal
+ t_b_777 peakVal 't_b_777+slope' baseVal
+ t_b_778 baseVal 't_b_778+slope' peakVal
+ t_b_779 peakVal 't_b_779+slope' baseVal
+ t_b_780 baseVal 't_b_780+slope' peakVal
+ t_b_781 peakVal 't_b_781+slope' baseVal
+ t_b_782 baseVal 't_b_782+slope' peakVal
+ t_b_783 peakVal 't_b_783+slope' baseVal
+ t_b_784 baseVal 't_b_784+slope' peakVal
+ t_b_785 peakVal 't_b_785+slope' baseVal
+ t_b_786 baseVal 't_b_786+slope' peakVal
+ t_b_787 peakVal 't_b_787+slope' baseVal
+ t_b_788 baseVal 't_b_788+slope' peakVal
+ t_b_789 peakVal 't_b_789+slope' baseVal
+ t_b_790 baseVal 't_b_790+slope' peakVal
+ t_b_791 peakVal 't_b_791+slope' baseVal
+ t_b_792 baseVal 't_b_792+slope' peakVal
+ t_b_793 peakVal 't_b_793+slope' baseVal
+ t_b_794 baseVal 't_b_794+slope' peakVal
+ t_b_795 peakVal 't_b_795+slope' baseVal
+ t_b_796 baseVal 't_b_796+slope' peakVal
+ t_b_797 peakVal 't_b_797+slope' baseVal
+ t_b_798 baseVal 't_b_798+slope' peakVal
+ t_b_799 peakVal 't_b_799+slope' baseVal




*circuit

XBUFFER_A Input_A A VDD VDD GND GND BUF_X8
XBUFFER_B Input_B B VDD VDD GND GND BUF_X8
XCGATE A B Z VDD VDD GND GND CGATE
XBUFFER_Z Z Output VDD VDD GND GND BUF_X8
C_TERM Output GND 0.0779pF

.PROBE TRAN V(A) V(B) V(Z)
.TRAN 0.1ps tend
.END
* circuit: cgate_test
simulator lang=spice

*.PARAM pw=<sed>pw<sed>as
.PARAM supp=0.8V slope=0.1fs
.PARAM t_init0=0.1ns t_init1=0.174ns
.PARAM baseVal=0V peakVal=0.8V tend=8100.0ns


.LIB /home/s11777724/involution_tool_library_files/backend/spice/fet.inc CMG

* main circuit
.INCLUDE /home/s11777724/involution_tool_library_files/backend/spice/cell/BUF_X8.sp
.INCLUDE cgate.sp

**** SPECTRE Back Annotation
.option spef='/home/s11777724/JS/idm_evaluation/cgate_test/place_and_route/cgate_test_restitch.spef'
****

.TEMP 25
.OPTION
+ INGOLD=2
+ PARHIER=LOCAL
*+ POST=CSDF
+ PROBE
+ BRIEF
+ ACCURATE
+ ABSVAR=0.0001
+ DVDT=2
+ RELTOL=1e-11
*+ DELMAX=100fs
+ dc_pivot_check=yes

* vdd
VDD VDD GND 0.8v

.PARAM t_a_0=10ns
.PARAM t_a_1=23.333333ns
.PARAM t_a_2=30ns
.PARAM t_a_3=43.333333ns
.PARAM t_a_4=50ns
.PARAM t_a_5=63.333333ns
.PARAM t_a_6=70ns
.PARAM t_a_7=83.333333ns
.PARAM t_a_8=90ns
.PARAM t_a_9=103.333333ns
.PARAM t_a_10=110ns
.PARAM t_a_11=123.333333ns
.PARAM t_a_12=130ns
.PARAM t_a_13=143.333333ns
.PARAM t_a_14=150ns
.PARAM t_a_15=163.333333ns
.PARAM t_a_16=170ns
.PARAM t_a_17=183.333333ns
.PARAM t_a_18=190ns
.PARAM t_a_19=203.333333ns
.PARAM t_a_20=210ns
.PARAM t_a_21=223.333333ns
.PARAM t_a_22=230ns
.PARAM t_a_23=243.333333ns
.PARAM t_a_24=250ns
.PARAM t_a_25=263.333333ns
.PARAM t_a_26=270ns
.PARAM t_a_27=283.333333ns
.PARAM t_a_28=290ns
.PARAM t_a_29=303.333333ns
.PARAM t_a_30=310ns
.PARAM t_a_31=323.333333ns
.PARAM t_a_32=330ns
.PARAM t_a_33=343.333333ns
.PARAM t_a_34=350ns
.PARAM t_a_35=363.333333ns
.PARAM t_a_36=370ns
.PARAM t_a_37=383.333333ns
.PARAM t_a_38=390ns
.PARAM t_a_39=403.333333ns
.PARAM t_a_40=410ns
.PARAM t_a_41=423.333333ns
.PARAM t_a_42=430ns
.PARAM t_a_43=443.333333ns
.PARAM t_a_44=450ns
.PARAM t_a_45=463.333333ns
.PARAM t_a_46=470ns
.PARAM t_a_47=483.333333ns
.PARAM t_a_48=490ns
.PARAM t_a_49=503.333333ns
.PARAM t_a_50=510ns
.PARAM t_a_51=523.333333ns
.PARAM t_a_52=530ns
.PARAM t_a_53=543.333333ns
.PARAM t_a_54=550ns
.PARAM t_a_55=563.333333ns
.PARAM t_a_56=570ns
.PARAM t_a_57=583.333333ns
.PARAM t_a_58=590ns
.PARAM t_a_59=603.333333ns
.PARAM t_a_60=610ns
.PARAM t_a_61=623.333333ns
.PARAM t_a_62=630ns
.PARAM t_a_63=643.333333ns
.PARAM t_a_64=650ns
.PARAM t_a_65=663.333333ns
.PARAM t_a_66=670ns
.PARAM t_a_67=683.333333ns
.PARAM t_a_68=690ns
.PARAM t_a_69=703.333333ns
.PARAM t_a_70=710ns
.PARAM t_a_71=723.333333ns
.PARAM t_a_72=730ns
.PARAM t_a_73=743.333333ns
.PARAM t_a_74=750ns
.PARAM t_a_75=763.333333ns
.PARAM t_a_76=770ns
.PARAM t_a_77=783.333333ns
.PARAM t_a_78=790ns
.PARAM t_a_79=803.333333ns
.PARAM t_a_80=810ns
.PARAM t_a_81=823.333333ns
.PARAM t_a_82=830ns
.PARAM t_a_83=843.333333ns
.PARAM t_a_84=850ns
.PARAM t_a_85=863.333333ns
.PARAM t_a_86=870ns
.PARAM t_a_87=883.333333ns
.PARAM t_a_88=890ns
.PARAM t_a_89=903.333333ns
.PARAM t_a_90=910ns
.PARAM t_a_91=923.333333ns
.PARAM t_a_92=930ns
.PARAM t_a_93=943.333333ns
.PARAM t_a_94=950ns
.PARAM t_a_95=963.333333ns
.PARAM t_a_96=970ns
.PARAM t_a_97=983.333333ns
.PARAM t_a_98=990ns
.PARAM t_a_99=1003.333333ns
.PARAM t_a_100=1010ns
.PARAM t_a_101=1023.333333ns
.PARAM t_a_102=1030ns
.PARAM t_a_103=1043.333333ns
.PARAM t_a_104=1050ns
.PARAM t_a_105=1063.333333ns
.PARAM t_a_106=1070ns
.PARAM t_a_107=1083.333333ns
.PARAM t_a_108=1090ns
.PARAM t_a_109=1103.333333ns
.PARAM t_a_110=1110ns
.PARAM t_a_111=1123.333333ns
.PARAM t_a_112=1130ns
.PARAM t_a_113=1143.333333ns
.PARAM t_a_114=1150ns
.PARAM t_a_115=1163.333333ns
.PARAM t_a_116=1170ns
.PARAM t_a_117=1183.333333ns
.PARAM t_a_118=1190ns
.PARAM t_a_119=1203.333333ns
.PARAM t_a_120=1210ns
.PARAM t_a_121=1223.333333ns
.PARAM t_a_122=1230ns
.PARAM t_a_123=1243.333333ns
.PARAM t_a_124=1250ns
.PARAM t_a_125=1263.333333ns
.PARAM t_a_126=1270ns
.PARAM t_a_127=1283.333333ns
.PARAM t_a_128=1290ns
.PARAM t_a_129=1303.333333ns
.PARAM t_a_130=1310ns
.PARAM t_a_131=1323.333333ns
.PARAM t_a_132=1330ns
.PARAM t_a_133=1343.333333ns
.PARAM t_a_134=1350ns
.PARAM t_a_135=1363.333333ns
.PARAM t_a_136=1370ns
.PARAM t_a_137=1383.333333ns
.PARAM t_a_138=1390ns
.PARAM t_a_139=1403.333333ns
.PARAM t_a_140=1410ns
.PARAM t_a_141=1423.333333ns
.PARAM t_a_142=1430ns
.PARAM t_a_143=1443.333333ns
.PARAM t_a_144=1450ns
.PARAM t_a_145=1463.333333ns
.PARAM t_a_146=1470ns
.PARAM t_a_147=1483.333333ns
.PARAM t_a_148=1490ns
.PARAM t_a_149=1503.333333ns
.PARAM t_a_150=1510ns
.PARAM t_a_151=1523.333333ns
.PARAM t_a_152=1530ns
.PARAM t_a_153=1543.333333ns
.PARAM t_a_154=1550ns
.PARAM t_a_155=1563.333333ns
.PARAM t_a_156=1570ns
.PARAM t_a_157=1583.333333ns
.PARAM t_a_158=1590ns
.PARAM t_a_159=1603.333333ns
.PARAM t_a_160=1610ns
.PARAM t_a_161=1623.333333ns
.PARAM t_a_162=1630ns
.PARAM t_a_163=1643.333333ns
.PARAM t_a_164=1650ns
.PARAM t_a_165=1663.333333ns
.PARAM t_a_166=1670ns
.PARAM t_a_167=1683.333333ns
.PARAM t_a_168=1690ns
.PARAM t_a_169=1703.333333ns
.PARAM t_a_170=1710ns
.PARAM t_a_171=1723.333333ns
.PARAM t_a_172=1730ns
.PARAM t_a_173=1743.333333ns
.PARAM t_a_174=1750ns
.PARAM t_a_175=1763.333333ns
.PARAM t_a_176=1770ns
.PARAM t_a_177=1783.333333ns
.PARAM t_a_178=1790ns
.PARAM t_a_179=1803.333333ns
.PARAM t_a_180=1810ns
.PARAM t_a_181=1823.333333ns
.PARAM t_a_182=1830ns
.PARAM t_a_183=1843.333333ns
.PARAM t_a_184=1850ns
.PARAM t_a_185=1863.333333ns
.PARAM t_a_186=1870ns
.PARAM t_a_187=1883.333333ns
.PARAM t_a_188=1890ns
.PARAM t_a_189=1903.333333ns
.PARAM t_a_190=1910ns
.PARAM t_a_191=1923.333333ns
.PARAM t_a_192=1930ns
.PARAM t_a_193=1943.333333ns
.PARAM t_a_194=1950ns
.PARAM t_a_195=1963.333333ns
.PARAM t_a_196=1970ns
.PARAM t_a_197=1983.333333ns
.PARAM t_a_198=1990ns
.PARAM t_a_199=2003.333333ns
.PARAM t_a_200=2010ns
.PARAM t_a_201=2023.333333ns
.PARAM t_a_202=2030ns
.PARAM t_a_203=2043.333333ns
.PARAM t_a_204=2050ns
.PARAM t_a_205=2063.333333ns
.PARAM t_a_206=2070ns
.PARAM t_a_207=2083.333333ns
.PARAM t_a_208=2090ns
.PARAM t_a_209=2103.333333ns
.PARAM t_a_210=2110ns
.PARAM t_a_211=2123.333333ns
.PARAM t_a_212=2130ns
.PARAM t_a_213=2143.333333ns
.PARAM t_a_214=2150ns
.PARAM t_a_215=2163.333333ns
.PARAM t_a_216=2170ns
.PARAM t_a_217=2183.333333ns
.PARAM t_a_218=2190ns
.PARAM t_a_219=2203.333333ns
.PARAM t_a_220=2210ns
.PARAM t_a_221=2223.333333ns
.PARAM t_a_222=2230ns
.PARAM t_a_223=2243.333333ns
.PARAM t_a_224=2250ns
.PARAM t_a_225=2263.333333ns
.PARAM t_a_226=2270ns
.PARAM t_a_227=2283.333333ns
.PARAM t_a_228=2290ns
.PARAM t_a_229=2303.333333ns
.PARAM t_a_230=2310ns
.PARAM t_a_231=2323.333333ns
.PARAM t_a_232=2330ns
.PARAM t_a_233=2343.333333ns
.PARAM t_a_234=2350ns
.PARAM t_a_235=2363.333333ns
.PARAM t_a_236=2370ns
.PARAM t_a_237=2383.333333ns
.PARAM t_a_238=2390ns
.PARAM t_a_239=2403.333333ns
.PARAM t_a_240=2410ns
.PARAM t_a_241=2423.333333ns
.PARAM t_a_242=2430ns
.PARAM t_a_243=2443.333333ns
.PARAM t_a_244=2450ns
.PARAM t_a_245=2463.333333ns
.PARAM t_a_246=2470ns
.PARAM t_a_247=2483.333333ns
.PARAM t_a_248=2490ns
.PARAM t_a_249=2503.333333ns
.PARAM t_a_250=2510ns
.PARAM t_a_251=2523.333333ns
.PARAM t_a_252=2530ns
.PARAM t_a_253=2543.333333ns
.PARAM t_a_254=2550ns
.PARAM t_a_255=2563.333333ns
.PARAM t_a_256=2570ns
.PARAM t_a_257=2583.333333ns
.PARAM t_a_258=2590ns
.PARAM t_a_259=2603.333333ns
.PARAM t_a_260=2610ns
.PARAM t_a_261=2623.333333ns
.PARAM t_a_262=2630ns
.PARAM t_a_263=2643.333333ns
.PARAM t_a_264=2650ns
.PARAM t_a_265=2663.333333ns
.PARAM t_a_266=2670ns
.PARAM t_a_267=2683.333333ns
.PARAM t_a_268=2690ns
.PARAM t_a_269=2703.333333ns
.PARAM t_a_270=2710ns
.PARAM t_a_271=2723.333333ns
.PARAM t_a_272=2730ns
.PARAM t_a_273=2743.333333ns
.PARAM t_a_274=2750ns
.PARAM t_a_275=2763.333333ns
.PARAM t_a_276=2770ns
.PARAM t_a_277=2783.333333ns
.PARAM t_a_278=2790ns
.PARAM t_a_279=2803.333333ns
.PARAM t_a_280=2810ns
.PARAM t_a_281=2823.333333ns
.PARAM t_a_282=2830ns
.PARAM t_a_283=2843.333333ns
.PARAM t_a_284=2850ns
.PARAM t_a_285=2863.333333ns
.PARAM t_a_286=2870ns
.PARAM t_a_287=2883.333333ns
.PARAM t_a_288=2890ns
.PARAM t_a_289=2903.333333ns
.PARAM t_a_290=2910ns
.PARAM t_a_291=2923.333333ns
.PARAM t_a_292=2930ns
.PARAM t_a_293=2943.333333ns
.PARAM t_a_294=2950ns
.PARAM t_a_295=2963.333333ns
.PARAM t_a_296=2970ns
.PARAM t_a_297=2983.333333ns
.PARAM t_a_298=2990ns
.PARAM t_a_299=3003.333333ns
.PARAM t_a_300=3010ns
.PARAM t_a_301=3023.333333ns
.PARAM t_a_302=3030ns
.PARAM t_a_303=3043.333333ns
.PARAM t_a_304=3050ns
.PARAM t_a_305=3063.333333ns
.PARAM t_a_306=3070ns
.PARAM t_a_307=3083.333333ns
.PARAM t_a_308=3090ns
.PARAM t_a_309=3103.333333ns
.PARAM t_a_310=3110ns
.PARAM t_a_311=3123.333333ns
.PARAM t_a_312=3130ns
.PARAM t_a_313=3143.333333ns
.PARAM t_a_314=3150ns
.PARAM t_a_315=3163.333333ns
.PARAM t_a_316=3170ns
.PARAM t_a_317=3183.333333ns
.PARAM t_a_318=3190ns
.PARAM t_a_319=3203.333333ns
.PARAM t_a_320=3210ns
.PARAM t_a_321=3223.333333ns
.PARAM t_a_322=3230ns
.PARAM t_a_323=3243.333333ns
.PARAM t_a_324=3250ns
.PARAM t_a_325=3263.333333ns
.PARAM t_a_326=3270ns
.PARAM t_a_327=3283.333333ns
.PARAM t_a_328=3290ns
.PARAM t_a_329=3303.333333ns
.PARAM t_a_330=3310ns
.PARAM t_a_331=3323.333333ns
.PARAM t_a_332=3330ns
.PARAM t_a_333=3343.333333ns
.PARAM t_a_334=3350ns
.PARAM t_a_335=3363.333333ns
.PARAM t_a_336=3370ns
.PARAM t_a_337=3383.333333ns
.PARAM t_a_338=3390ns
.PARAM t_a_339=3403.333333ns
.PARAM t_a_340=3410ns
.PARAM t_a_341=3423.333333ns
.PARAM t_a_342=3430ns
.PARAM t_a_343=3443.333333ns
.PARAM t_a_344=3450ns
.PARAM t_a_345=3463.333333ns
.PARAM t_a_346=3470ns
.PARAM t_a_347=3483.333333ns
.PARAM t_a_348=3490ns
.PARAM t_a_349=3503.333333ns
.PARAM t_a_350=3510ns
.PARAM t_a_351=3523.333333ns
.PARAM t_a_352=3530ns
.PARAM t_a_353=3543.333333ns
.PARAM t_a_354=3550ns
.PARAM t_a_355=3563.333333ns
.PARAM t_a_356=3570ns
.PARAM t_a_357=3583.333333ns
.PARAM t_a_358=3590ns
.PARAM t_a_359=3603.333333ns
.PARAM t_a_360=3610ns
.PARAM t_a_361=3623.333333ns
.PARAM t_a_362=3630ns
.PARAM t_a_363=3643.333333ns
.PARAM t_a_364=3650ns
.PARAM t_a_365=3663.333333ns
.PARAM t_a_366=3670ns
.PARAM t_a_367=3683.333333ns
.PARAM t_a_368=3690ns
.PARAM t_a_369=3703.333333ns
.PARAM t_a_370=3710ns
.PARAM t_a_371=3723.333333ns
.PARAM t_a_372=3730ns
.PARAM t_a_373=3743.333333ns
.PARAM t_a_374=3750ns
.PARAM t_a_375=3763.333333ns
.PARAM t_a_376=3770ns
.PARAM t_a_377=3783.333333ns
.PARAM t_a_378=3790ns
.PARAM t_a_379=3803.333333ns
.PARAM t_a_380=3810ns
.PARAM t_a_381=3823.333333ns
.PARAM t_a_382=3830ns
.PARAM t_a_383=3843.333333ns
.PARAM t_a_384=3850ns
.PARAM t_a_385=3863.333333ns
.PARAM t_a_386=3870ns
.PARAM t_a_387=3883.333333ns
.PARAM t_a_388=3890ns
.PARAM t_a_389=3903.333333ns
.PARAM t_a_390=3910ns
.PARAM t_a_391=3923.333333ns
.PARAM t_a_392=3930ns
.PARAM t_a_393=3943.333333ns
.PARAM t_a_394=3950ns
.PARAM t_a_395=3963.333333ns
.PARAM t_a_396=3970ns
.PARAM t_a_397=3983.333333ns
.PARAM t_a_398=3990ns
.PARAM t_a_399=4003.333333ns
.PARAM t_a_400=4010ns
.PARAM t_a_401=4023.333333ns
.PARAM t_a_402=4030ns
.PARAM t_a_403=4043.333333ns
.PARAM t_a_404=4050ns
.PARAM t_a_405=4063.333333ns
.PARAM t_a_406=4070ns
.PARAM t_a_407=4083.333333ns
.PARAM t_a_408=4090ns
.PARAM t_a_409=4103.333333ns
.PARAM t_a_410=4110ns
.PARAM t_a_411=4123.333333ns
.PARAM t_a_412=4130ns
.PARAM t_a_413=4143.333333ns
.PARAM t_a_414=4150ns
.PARAM t_a_415=4163.333333ns
.PARAM t_a_416=4170ns
.PARAM t_a_417=4183.333333ns
.PARAM t_a_418=4190ns
.PARAM t_a_419=4203.333333ns
.PARAM t_a_420=4210ns
.PARAM t_a_421=4223.333333ns
.PARAM t_a_422=4230ns
.PARAM t_a_423=4243.333333ns
.PARAM t_a_424=4250ns
.PARAM t_a_425=4263.333333ns
.PARAM t_a_426=4270ns
.PARAM t_a_427=4283.333333ns
.PARAM t_a_428=4290ns
.PARAM t_a_429=4303.333333ns
.PARAM t_a_430=4310ns
.PARAM t_a_431=4323.333333ns
.PARAM t_a_432=4330ns
.PARAM t_a_433=4343.333333ns
.PARAM t_a_434=4350ns
.PARAM t_a_435=4363.333333ns
.PARAM t_a_436=4370ns
.PARAM t_a_437=4383.333333ns
.PARAM t_a_438=4390ns
.PARAM t_a_439=4403.333333ns
.PARAM t_a_440=4410ns
.PARAM t_a_441=4423.333333ns
.PARAM t_a_442=4430ns
.PARAM t_a_443=4443.333333ns
.PARAM t_a_444=4450ns
.PARAM t_a_445=4463.333333ns
.PARAM t_a_446=4470ns
.PARAM t_a_447=4483.333333ns
.PARAM t_a_448=4490ns
.PARAM t_a_449=4503.333333ns
.PARAM t_a_450=4510ns
.PARAM t_a_451=4523.333333ns
.PARAM t_a_452=4530ns
.PARAM t_a_453=4543.333333ns
.PARAM t_a_454=4550ns
.PARAM t_a_455=4563.333333ns
.PARAM t_a_456=4570ns
.PARAM t_a_457=4583.333333ns
.PARAM t_a_458=4590ns
.PARAM t_a_459=4603.333333ns
.PARAM t_a_460=4610ns
.PARAM t_a_461=4623.333333ns
.PARAM t_a_462=4630ns
.PARAM t_a_463=4643.333333ns
.PARAM t_a_464=4650ns
.PARAM t_a_465=4663.333333ns
.PARAM t_a_466=4670ns
.PARAM t_a_467=4683.333333ns
.PARAM t_a_468=4690ns
.PARAM t_a_469=4703.333333ns
.PARAM t_a_470=4710ns
.PARAM t_a_471=4723.333333ns
.PARAM t_a_472=4730ns
.PARAM t_a_473=4743.333333ns
.PARAM t_a_474=4750ns
.PARAM t_a_475=4763.333333ns
.PARAM t_a_476=4770ns
.PARAM t_a_477=4783.333333ns
.PARAM t_a_478=4790ns
.PARAM t_a_479=4803.333333ns
.PARAM t_a_480=4810ns
.PARAM t_a_481=4823.333333ns
.PARAM t_a_482=4830ns
.PARAM t_a_483=4843.333333ns
.PARAM t_a_484=4850ns
.PARAM t_a_485=4863.333333ns
.PARAM t_a_486=4870ns
.PARAM t_a_487=4883.333333ns
.PARAM t_a_488=4890ns
.PARAM t_a_489=4903.333333ns
.PARAM t_a_490=4910ns
.PARAM t_a_491=4923.333333ns
.PARAM t_a_492=4930ns
.PARAM t_a_493=4943.333333ns
.PARAM t_a_494=4950ns
.PARAM t_a_495=4963.333333ns
.PARAM t_a_496=4970ns
.PARAM t_a_497=4983.333333ns
.PARAM t_a_498=4990ns
.PARAM t_a_499=5003.333333ns
.PARAM t_a_500=5010ns
.PARAM t_a_501=5023.333333ns
.PARAM t_a_502=5030ns
.PARAM t_a_503=5043.333333ns
.PARAM t_a_504=5050ns
.PARAM t_a_505=5063.333333ns
.PARAM t_a_506=5070ns
.PARAM t_a_507=5083.333333ns
.PARAM t_a_508=5090ns
.PARAM t_a_509=5103.333333ns
.PARAM t_a_510=5110ns
.PARAM t_a_511=5123.333333ns
.PARAM t_a_512=5130ns
.PARAM t_a_513=5143.333333ns
.PARAM t_a_514=5150ns
.PARAM t_a_515=5163.333333ns
.PARAM t_a_516=5170ns
.PARAM t_a_517=5183.333333ns
.PARAM t_a_518=5190ns
.PARAM t_a_519=5203.333333ns
.PARAM t_a_520=5210ns
.PARAM t_a_521=5223.333333ns
.PARAM t_a_522=5230ns
.PARAM t_a_523=5243.333333ns
.PARAM t_a_524=5250ns
.PARAM t_a_525=5263.333333ns
.PARAM t_a_526=5270ns
.PARAM t_a_527=5283.333333ns
.PARAM t_a_528=5290ns
.PARAM t_a_529=5303.333333ns
.PARAM t_a_530=5310ns
.PARAM t_a_531=5323.333333ns
.PARAM t_a_532=5330ns
.PARAM t_a_533=5343.333333ns
.PARAM t_a_534=5350ns
.PARAM t_a_535=5363.333333ns
.PARAM t_a_536=5370ns
.PARAM t_a_537=5383.333333ns
.PARAM t_a_538=5390ns
.PARAM t_a_539=5403.333333ns
.PARAM t_a_540=5410ns
.PARAM t_a_541=5423.333333ns
.PARAM t_a_542=5430ns
.PARAM t_a_543=5443.333333ns
.PARAM t_a_544=5450ns
.PARAM t_a_545=5463.333333ns
.PARAM t_a_546=5470ns
.PARAM t_a_547=5483.333333ns
.PARAM t_a_548=5490ns
.PARAM t_a_549=5503.333333ns
.PARAM t_a_550=5510ns
.PARAM t_a_551=5523.333333ns
.PARAM t_a_552=5530ns
.PARAM t_a_553=5543.333333ns
.PARAM t_a_554=5550ns
.PARAM t_a_555=5563.333333ns
.PARAM t_a_556=5570ns
.PARAM t_a_557=5583.333333ns
.PARAM t_a_558=5590ns
.PARAM t_a_559=5603.333333ns
.PARAM t_a_560=5610ns
.PARAM t_a_561=5623.333333ns
.PARAM t_a_562=5630ns
.PARAM t_a_563=5643.333333ns
.PARAM t_a_564=5650ns
.PARAM t_a_565=5663.333333ns
.PARAM t_a_566=5670ns
.PARAM t_a_567=5683.333333ns
.PARAM t_a_568=5690ns
.PARAM t_a_569=5703.333333ns
.PARAM t_a_570=5710ns
.PARAM t_a_571=5723.333333ns
.PARAM t_a_572=5730ns
.PARAM t_a_573=5743.333333ns
.PARAM t_a_574=5750ns
.PARAM t_a_575=5763.333333ns
.PARAM t_a_576=5770ns
.PARAM t_a_577=5783.333333ns
.PARAM t_a_578=5790ns
.PARAM t_a_579=5803.333333ns
.PARAM t_a_580=5810ns
.PARAM t_a_581=5823.333333ns
.PARAM t_a_582=5830ns
.PARAM t_a_583=5843.333333ns
.PARAM t_a_584=5850ns
.PARAM t_a_585=5863.333333ns
.PARAM t_a_586=5870ns
.PARAM t_a_587=5883.333333ns
.PARAM t_a_588=5890ns
.PARAM t_a_589=5903.333333ns
.PARAM t_a_590=5910ns
.PARAM t_a_591=5923.333333ns
.PARAM t_a_592=5930ns
.PARAM t_a_593=5943.333333ns
.PARAM t_a_594=5950ns
.PARAM t_a_595=5963.333333ns
.PARAM t_a_596=5970ns
.PARAM t_a_597=5983.333333ns
.PARAM t_a_598=5990ns
.PARAM t_a_599=6003.333333ns
.PARAM t_a_600=6010ns
.PARAM t_a_601=6023.333333ns
.PARAM t_a_602=6030ns
.PARAM t_a_603=6043.333333ns
.PARAM t_a_604=6050ns
.PARAM t_a_605=6063.333333ns
.PARAM t_a_606=6070ns
.PARAM t_a_607=6083.333333ns
.PARAM t_a_608=6090ns
.PARAM t_a_609=6103.333333ns
.PARAM t_a_610=6110ns
.PARAM t_a_611=6123.333333ns
.PARAM t_a_612=6130ns
.PARAM t_a_613=6143.333333ns
.PARAM t_a_614=6150ns
.PARAM t_a_615=6163.333333ns
.PARAM t_a_616=6170ns
.PARAM t_a_617=6183.333333ns
.PARAM t_a_618=6190ns
.PARAM t_a_619=6203.333333ns
.PARAM t_a_620=6210ns
.PARAM t_a_621=6223.333333ns
.PARAM t_a_622=6230ns
.PARAM t_a_623=6243.333333ns
.PARAM t_a_624=6250ns
.PARAM t_a_625=6263.333333ns
.PARAM t_a_626=6270ns
.PARAM t_a_627=6283.333333ns
.PARAM t_a_628=6290ns
.PARAM t_a_629=6303.333333ns
.PARAM t_a_630=6310ns
.PARAM t_a_631=6323.333333ns
.PARAM t_a_632=6330ns
.PARAM t_a_633=6343.333333ns
.PARAM t_a_634=6350ns
.PARAM t_a_635=6363.333333ns
.PARAM t_a_636=6370ns
.PARAM t_a_637=6383.333333ns
.PARAM t_a_638=6390ns
.PARAM t_a_639=6403.333333ns
.PARAM t_a_640=6410ns
.PARAM t_a_641=6423.333333ns
.PARAM t_a_642=6430ns
.PARAM t_a_643=6443.333333ns
.PARAM t_a_644=6450ns
.PARAM t_a_645=6463.333333ns
.PARAM t_a_646=6470ns
.PARAM t_a_647=6483.333333ns
.PARAM t_a_648=6490ns
.PARAM t_a_649=6503.333333ns
.PARAM t_a_650=6510ns
.PARAM t_a_651=6523.333333ns
.PARAM t_a_652=6530ns
.PARAM t_a_653=6543.333333ns
.PARAM t_a_654=6550ns
.PARAM t_a_655=6563.333333ns
.PARAM t_a_656=6570ns
.PARAM t_a_657=6583.333333ns
.PARAM t_a_658=6590ns
.PARAM t_a_659=6603.333333ns
.PARAM t_a_660=6610ns
.PARAM t_a_661=6623.333333ns
.PARAM t_a_662=6630ns
.PARAM t_a_663=6643.333333ns
.PARAM t_a_664=6650ns
.PARAM t_a_665=6663.333333ns
.PARAM t_a_666=6670ns
.PARAM t_a_667=6683.333333ns
.PARAM t_a_668=6690ns
.PARAM t_a_669=6703.333333ns
.PARAM t_a_670=6710ns
.PARAM t_a_671=6723.333333ns
.PARAM t_a_672=6730ns
.PARAM t_a_673=6743.333333ns
.PARAM t_a_674=6750ns
.PARAM t_a_675=6763.333333ns
.PARAM t_a_676=6770ns
.PARAM t_a_677=6783.333333ns
.PARAM t_a_678=6790ns
.PARAM t_a_679=6803.333333ns
.PARAM t_a_680=6810ns
.PARAM t_a_681=6823.333333ns
.PARAM t_a_682=6830ns
.PARAM t_a_683=6843.333333ns
.PARAM t_a_684=6850ns
.PARAM t_a_685=6863.333333ns
.PARAM t_a_686=6870ns
.PARAM t_a_687=6883.333333ns
.PARAM t_a_688=6890ns
.PARAM t_a_689=6903.333333ns
.PARAM t_a_690=6910ns
.PARAM t_a_691=6923.333333ns
.PARAM t_a_692=6930ns
.PARAM t_a_693=6943.333333ns
.PARAM t_a_694=6950ns
.PARAM t_a_695=6963.333333ns
.PARAM t_a_696=6970ns
.PARAM t_a_697=6983.333333ns
.PARAM t_a_698=6990ns
.PARAM t_a_699=7003.333333ns
.PARAM t_a_700=7010ns
.PARAM t_a_701=7023.333333ns
.PARAM t_a_702=7030ns
.PARAM t_a_703=7043.333333ns
.PARAM t_a_704=7050ns
.PARAM t_a_705=7063.333333ns
.PARAM t_a_706=7070ns
.PARAM t_a_707=7083.333333ns
.PARAM t_a_708=7090ns
.PARAM t_a_709=7103.333333ns
.PARAM t_a_710=7110ns
.PARAM t_a_711=7123.333333ns
.PARAM t_a_712=7130ns
.PARAM t_a_713=7143.333333ns
.PARAM t_a_714=7150ns
.PARAM t_a_715=7163.333333ns
.PARAM t_a_716=7170ns
.PARAM t_a_717=7183.333333ns
.PARAM t_a_718=7190ns
.PARAM t_a_719=7203.333333ns
.PARAM t_a_720=7210ns
.PARAM t_a_721=7223.333333ns
.PARAM t_a_722=7230ns
.PARAM t_a_723=7243.333333ns
.PARAM t_a_724=7250ns
.PARAM t_a_725=7263.333333ns
.PARAM t_a_726=7270ns
.PARAM t_a_727=7283.333333ns
.PARAM t_a_728=7290ns
.PARAM t_a_729=7303.333333ns
.PARAM t_a_730=7310ns
.PARAM t_a_731=7323.333333ns
.PARAM t_a_732=7330ns
.PARAM t_a_733=7343.333333ns
.PARAM t_a_734=7350ns
.PARAM t_a_735=7363.333333ns
.PARAM t_a_736=7370ns
.PARAM t_a_737=7383.333333ns
.PARAM t_a_738=7390ns
.PARAM t_a_739=7403.333333ns
.PARAM t_a_740=7410ns
.PARAM t_a_741=7423.333333ns
.PARAM t_a_742=7430ns
.PARAM t_a_743=7443.333333ns
.PARAM t_a_744=7450ns
.PARAM t_a_745=7463.333333ns
.PARAM t_a_746=7470ns
.PARAM t_a_747=7483.333333ns
.PARAM t_a_748=7490ns
.PARAM t_a_749=7503.333333ns
.PARAM t_a_750=7510ns
.PARAM t_a_751=7523.333333ns
.PARAM t_a_752=7530ns
.PARAM t_a_753=7543.333333ns
.PARAM t_a_754=7550ns
.PARAM t_a_755=7563.333333ns
.PARAM t_a_756=7570ns
.PARAM t_a_757=7583.333333ns
.PARAM t_a_758=7590ns
.PARAM t_a_759=7603.333333ns
.PARAM t_a_760=7610ns
.PARAM t_a_761=7623.333333ns
.PARAM t_a_762=7630ns
.PARAM t_a_763=7643.333333ns
.PARAM t_a_764=7650ns
.PARAM t_a_765=7663.333333ns
.PARAM t_a_766=7670ns
.PARAM t_a_767=7683.333333ns
.PARAM t_a_768=7690ns
.PARAM t_a_769=7703.333333ns
.PARAM t_a_770=7710ns
.PARAM t_a_771=7723.333333ns
.PARAM t_a_772=7730ns
.PARAM t_a_773=7743.333333ns
.PARAM t_a_774=7750ns
.PARAM t_a_775=7763.333333ns
.PARAM t_a_776=7770ns
.PARAM t_a_777=7783.333333ns
.PARAM t_a_778=7790ns
.PARAM t_a_779=7803.333333ns
.PARAM t_a_780=7810ns
.PARAM t_a_781=7823.333333ns
.PARAM t_a_782=7830ns
.PARAM t_a_783=7843.333333ns
.PARAM t_a_784=7850ns
.PARAM t_a_785=7863.333333ns
.PARAM t_a_786=7870ns
.PARAM t_a_787=7883.333333ns
.PARAM t_a_788=7890ns
.PARAM t_a_789=7903.333333ns
.PARAM t_a_790=7910ns
.PARAM t_a_791=7923.333333ns
.PARAM t_a_792=7930ns
.PARAM t_a_793=7943.333333ns
.PARAM t_a_794=7950ns
.PARAM t_a_795=7963.333333ns
.PARAM t_a_796=7970ns
.PARAM t_a_797=7983.333333ns
.PARAM t_a_798=7990ns
.PARAM t_a_799=8003.333333ns
.PARAM t_b_0=9.8ns
.PARAM t_b_1=16.666667ns
.PARAM t_b_2=29.801ns
.PARAM t_b_3=36.666667ns
.PARAM t_b_4=49.802ns
.PARAM t_b_5=56.666667ns
.PARAM t_b_6=69.803ns
.PARAM t_b_7=76.666667ns
.PARAM t_b_8=89.804ns
.PARAM t_b_9=96.666667ns
.PARAM t_b_10=109.805ns
.PARAM t_b_11=116.666667ns
.PARAM t_b_12=129.806ns
.PARAM t_b_13=136.666667ns
.PARAM t_b_14=149.807ns
.PARAM t_b_15=156.666667ns
.PARAM t_b_16=169.808ns
.PARAM t_b_17=176.666667ns
.PARAM t_b_18=189.809ns
.PARAM t_b_19=196.666667ns
.PARAM t_b_20=209.81ns
.PARAM t_b_21=216.666667ns
.PARAM t_b_22=229.811ns
.PARAM t_b_23=236.666667ns
.PARAM t_b_24=249.812ns
.PARAM t_b_25=256.666667ns
.PARAM t_b_26=269.813ns
.PARAM t_b_27=276.666667ns
.PARAM t_b_28=289.814ns
.PARAM t_b_29=296.666667ns
.PARAM t_b_30=309.815ns
.PARAM t_b_31=316.666667ns
.PARAM t_b_32=329.816ns
.PARAM t_b_33=336.666667ns
.PARAM t_b_34=349.817ns
.PARAM t_b_35=356.666667ns
.PARAM t_b_36=369.818ns
.PARAM t_b_37=376.666667ns
.PARAM t_b_38=389.819ns
.PARAM t_b_39=396.666667ns
.PARAM t_b_40=409.82ns
.PARAM t_b_41=416.666667ns
.PARAM t_b_42=429.821ns
.PARAM t_b_43=436.666667ns
.PARAM t_b_44=449.822ns
.PARAM t_b_45=456.666667ns
.PARAM t_b_46=469.823ns
.PARAM t_b_47=476.666667ns
.PARAM t_b_48=489.824ns
.PARAM t_b_49=496.666667ns
.PARAM t_b_50=509.825ns
.PARAM t_b_51=516.666667ns
.PARAM t_b_52=529.826ns
.PARAM t_b_53=536.666667ns
.PARAM t_b_54=549.827ns
.PARAM t_b_55=556.666667ns
.PARAM t_b_56=569.828ns
.PARAM t_b_57=576.666667ns
.PARAM t_b_58=589.829ns
.PARAM t_b_59=596.666667ns
.PARAM t_b_60=609.83ns
.PARAM t_b_61=616.666667ns
.PARAM t_b_62=629.831ns
.PARAM t_b_63=636.666667ns
.PARAM t_b_64=649.832ns
.PARAM t_b_65=656.666667ns
.PARAM t_b_66=669.833ns
.PARAM t_b_67=676.666667ns
.PARAM t_b_68=689.834ns
.PARAM t_b_69=696.666667ns
.PARAM t_b_70=709.835ns
.PARAM t_b_71=716.666667ns
.PARAM t_b_72=729.836ns
.PARAM t_b_73=736.666667ns
.PARAM t_b_74=749.837ns
.PARAM t_b_75=756.666667ns
.PARAM t_b_76=769.838ns
.PARAM t_b_77=776.666667ns
.PARAM t_b_78=789.839ns
.PARAM t_b_79=796.666667ns
.PARAM t_b_80=809.84ns
.PARAM t_b_81=816.666667ns
.PARAM t_b_82=829.841ns
.PARAM t_b_83=836.666667ns
.PARAM t_b_84=849.842ns
.PARAM t_b_85=856.666667ns
.PARAM t_b_86=869.843ns
.PARAM t_b_87=876.666667ns
.PARAM t_b_88=889.844ns
.PARAM t_b_89=896.666667ns
.PARAM t_b_90=909.845ns
.PARAM t_b_91=916.666667ns
.PARAM t_b_92=929.846ns
.PARAM t_b_93=936.666667ns
.PARAM t_b_94=949.847ns
.PARAM t_b_95=956.666667ns
.PARAM t_b_96=969.848ns
.PARAM t_b_97=976.666667ns
.PARAM t_b_98=989.849ns
.PARAM t_b_99=996.666667ns
.PARAM t_b_100=1009.85ns
.PARAM t_b_101=1016.666667ns
.PARAM t_b_102=1029.851ns
.PARAM t_b_103=1036.666667ns
.PARAM t_b_104=1049.852ns
.PARAM t_b_105=1056.666667ns
.PARAM t_b_106=1069.853ns
.PARAM t_b_107=1076.666667ns
.PARAM t_b_108=1089.854ns
.PARAM t_b_109=1096.666667ns
.PARAM t_b_110=1109.855ns
.PARAM t_b_111=1116.666667ns
.PARAM t_b_112=1129.856ns
.PARAM t_b_113=1136.666667ns
.PARAM t_b_114=1149.857ns
.PARAM t_b_115=1156.666667ns
.PARAM t_b_116=1169.858ns
.PARAM t_b_117=1176.666667ns
.PARAM t_b_118=1189.859ns
.PARAM t_b_119=1196.666667ns
.PARAM t_b_120=1209.86ns
.PARAM t_b_121=1216.666667ns
.PARAM t_b_122=1229.861ns
.PARAM t_b_123=1236.666667ns
.PARAM t_b_124=1249.862ns
.PARAM t_b_125=1256.666667ns
.PARAM t_b_126=1269.863ns
.PARAM t_b_127=1276.666667ns
.PARAM t_b_128=1289.864ns
.PARAM t_b_129=1296.666667ns
.PARAM t_b_130=1309.865ns
.PARAM t_b_131=1316.666667ns
.PARAM t_b_132=1329.866ns
.PARAM t_b_133=1336.666667ns
.PARAM t_b_134=1349.867ns
.PARAM t_b_135=1356.666667ns
.PARAM t_b_136=1369.868ns
.PARAM t_b_137=1376.666667ns
.PARAM t_b_138=1389.869ns
.PARAM t_b_139=1396.666667ns
.PARAM t_b_140=1409.87ns
.PARAM t_b_141=1416.666667ns
.PARAM t_b_142=1429.871ns
.PARAM t_b_143=1436.666667ns
.PARAM t_b_144=1449.872ns
.PARAM t_b_145=1456.666667ns
.PARAM t_b_146=1469.873ns
.PARAM t_b_147=1476.666667ns
.PARAM t_b_148=1489.874ns
.PARAM t_b_149=1496.666667ns
.PARAM t_b_150=1509.875ns
.PARAM t_b_151=1516.666667ns
.PARAM t_b_152=1529.876ns
.PARAM t_b_153=1536.666667ns
.PARAM t_b_154=1549.877ns
.PARAM t_b_155=1556.666667ns
.PARAM t_b_156=1569.878ns
.PARAM t_b_157=1576.666667ns
.PARAM t_b_158=1589.879ns
.PARAM t_b_159=1596.666667ns
.PARAM t_b_160=1609.88ns
.PARAM t_b_161=1616.666667ns
.PARAM t_b_162=1629.881ns
.PARAM t_b_163=1636.666667ns
.PARAM t_b_164=1649.882ns
.PARAM t_b_165=1656.666667ns
.PARAM t_b_166=1669.883ns
.PARAM t_b_167=1676.666667ns
.PARAM t_b_168=1689.884ns
.PARAM t_b_169=1696.666667ns
.PARAM t_b_170=1709.885ns
.PARAM t_b_171=1716.666667ns
.PARAM t_b_172=1729.886ns
.PARAM t_b_173=1736.666667ns
.PARAM t_b_174=1749.887ns
.PARAM t_b_175=1756.666667ns
.PARAM t_b_176=1769.888ns
.PARAM t_b_177=1776.666667ns
.PARAM t_b_178=1789.889ns
.PARAM t_b_179=1796.666667ns
.PARAM t_b_180=1809.89ns
.PARAM t_b_181=1816.666667ns
.PARAM t_b_182=1829.891ns
.PARAM t_b_183=1836.666667ns
.PARAM t_b_184=1849.892ns
.PARAM t_b_185=1856.666667ns
.PARAM t_b_186=1869.893ns
.PARAM t_b_187=1876.666667ns
.PARAM t_b_188=1889.894ns
.PARAM t_b_189=1896.666667ns
.PARAM t_b_190=1909.895ns
.PARAM t_b_191=1916.666667ns
.PARAM t_b_192=1929.896ns
.PARAM t_b_193=1936.666667ns
.PARAM t_b_194=1949.897ns
.PARAM t_b_195=1956.666667ns
.PARAM t_b_196=1969.898ns
.PARAM t_b_197=1976.666667ns
.PARAM t_b_198=1989.899ns
.PARAM t_b_199=1996.666667ns
.PARAM t_b_200=2009.9ns
.PARAM t_b_201=2016.666667ns
.PARAM t_b_202=2029.901ns
.PARAM t_b_203=2036.666667ns
.PARAM t_b_204=2049.902ns
.PARAM t_b_205=2056.666667ns
.PARAM t_b_206=2069.903ns
.PARAM t_b_207=2076.666667ns
.PARAM t_b_208=2089.904ns
.PARAM t_b_209=2096.666667ns
.PARAM t_b_210=2109.905ns
.PARAM t_b_211=2116.666667ns
.PARAM t_b_212=2129.906ns
.PARAM t_b_213=2136.666667ns
.PARAM t_b_214=2149.907ns
.PARAM t_b_215=2156.666667ns
.PARAM t_b_216=2169.908ns
.PARAM t_b_217=2176.666667ns
.PARAM t_b_218=2189.909ns
.PARAM t_b_219=2196.666667ns
.PARAM t_b_220=2209.91ns
.PARAM t_b_221=2216.666667ns
.PARAM t_b_222=2229.911ns
.PARAM t_b_223=2236.666667ns
.PARAM t_b_224=2249.912ns
.PARAM t_b_225=2256.666667ns
.PARAM t_b_226=2269.913ns
.PARAM t_b_227=2276.666667ns
.PARAM t_b_228=2289.914ns
.PARAM t_b_229=2296.666667ns
.PARAM t_b_230=2309.915ns
.PARAM t_b_231=2316.666667ns
.PARAM t_b_232=2329.916ns
.PARAM t_b_233=2336.666667ns
.PARAM t_b_234=2349.917ns
.PARAM t_b_235=2356.666667ns
.PARAM t_b_236=2369.918ns
.PARAM t_b_237=2376.666667ns
.PARAM t_b_238=2389.919ns
.PARAM t_b_239=2396.666667ns
.PARAM t_b_240=2409.92ns
.PARAM t_b_241=2416.666667ns
.PARAM t_b_242=2429.921ns
.PARAM t_b_243=2436.666667ns
.PARAM t_b_244=2449.922ns
.PARAM t_b_245=2456.666667ns
.PARAM t_b_246=2469.923ns
.PARAM t_b_247=2476.666667ns
.PARAM t_b_248=2489.924ns
.PARAM t_b_249=2496.666667ns
.PARAM t_b_250=2509.925ns
.PARAM t_b_251=2516.666667ns
.PARAM t_b_252=2529.926ns
.PARAM t_b_253=2536.666667ns
.PARAM t_b_254=2549.927ns
.PARAM t_b_255=2556.666667ns
.PARAM t_b_256=2569.928ns
.PARAM t_b_257=2576.666667ns
.PARAM t_b_258=2589.929ns
.PARAM t_b_259=2596.666667ns
.PARAM t_b_260=2609.93ns
.PARAM t_b_261=2616.666667ns
.PARAM t_b_262=2629.931ns
.PARAM t_b_263=2636.666667ns
.PARAM t_b_264=2649.932ns
.PARAM t_b_265=2656.666667ns
.PARAM t_b_266=2669.933ns
.PARAM t_b_267=2676.666667ns
.PARAM t_b_268=2689.934ns
.PARAM t_b_269=2696.666667ns
.PARAM t_b_270=2709.935ns
.PARAM t_b_271=2716.666667ns
.PARAM t_b_272=2729.936ns
.PARAM t_b_273=2736.666667ns
.PARAM t_b_274=2749.937ns
.PARAM t_b_275=2756.666667ns
.PARAM t_b_276=2769.938ns
.PARAM t_b_277=2776.666667ns
.PARAM t_b_278=2789.939ns
.PARAM t_b_279=2796.666667ns
.PARAM t_b_280=2809.94ns
.PARAM t_b_281=2816.666667ns
.PARAM t_b_282=2829.941ns
.PARAM t_b_283=2836.666667ns
.PARAM t_b_284=2849.942ns
.PARAM t_b_285=2856.666667ns
.PARAM t_b_286=2869.943ns
.PARAM t_b_287=2876.666667ns
.PARAM t_b_288=2889.944ns
.PARAM t_b_289=2896.666667ns
.PARAM t_b_290=2909.945ns
.PARAM t_b_291=2916.666667ns
.PARAM t_b_292=2929.946ns
.PARAM t_b_293=2936.666667ns
.PARAM t_b_294=2949.947ns
.PARAM t_b_295=2956.666667ns
.PARAM t_b_296=2969.948ns
.PARAM t_b_297=2976.666667ns
.PARAM t_b_298=2989.949ns
.PARAM t_b_299=2996.666667ns
.PARAM t_b_300=3009.95ns
.PARAM t_b_301=3016.666667ns
.PARAM t_b_302=3029.951ns
.PARAM t_b_303=3036.666667ns
.PARAM t_b_304=3049.952ns
.PARAM t_b_305=3056.666667ns
.PARAM t_b_306=3069.953ns
.PARAM t_b_307=3076.666667ns
.PARAM t_b_308=3089.954ns
.PARAM t_b_309=3096.666667ns
.PARAM t_b_310=3109.955ns
.PARAM t_b_311=3116.666667ns
.PARAM t_b_312=3129.956ns
.PARAM t_b_313=3136.666667ns
.PARAM t_b_314=3149.957ns
.PARAM t_b_315=3156.666667ns
.PARAM t_b_316=3169.958ns
.PARAM t_b_317=3176.666667ns
.PARAM t_b_318=3189.959ns
.PARAM t_b_319=3196.666667ns
.PARAM t_b_320=3209.96ns
.PARAM t_b_321=3216.666667ns
.PARAM t_b_322=3229.961ns
.PARAM t_b_323=3236.666667ns
.PARAM t_b_324=3249.962ns
.PARAM t_b_325=3256.666667ns
.PARAM t_b_326=3269.963ns
.PARAM t_b_327=3276.666667ns
.PARAM t_b_328=3289.964ns
.PARAM t_b_329=3296.666667ns
.PARAM t_b_330=3309.965ns
.PARAM t_b_331=3316.666667ns
.PARAM t_b_332=3329.966ns
.PARAM t_b_333=3336.666667ns
.PARAM t_b_334=3349.967ns
.PARAM t_b_335=3356.666667ns
.PARAM t_b_336=3369.968ns
.PARAM t_b_337=3376.666667ns
.PARAM t_b_338=3389.969ns
.PARAM t_b_339=3396.666667ns
.PARAM t_b_340=3409.97ns
.PARAM t_b_341=3416.666667ns
.PARAM t_b_342=3429.971ns
.PARAM t_b_343=3436.666667ns
.PARAM t_b_344=3449.972ns
.PARAM t_b_345=3456.666667ns
.PARAM t_b_346=3469.973ns
.PARAM t_b_347=3476.666667ns
.PARAM t_b_348=3489.974ns
.PARAM t_b_349=3496.666667ns
.PARAM t_b_350=3509.975ns
.PARAM t_b_351=3516.666667ns
.PARAM t_b_352=3529.976ns
.PARAM t_b_353=3536.666667ns
.PARAM t_b_354=3549.977ns
.PARAM t_b_355=3556.666667ns
.PARAM t_b_356=3569.978ns
.PARAM t_b_357=3576.666667ns
.PARAM t_b_358=3589.979ns
.PARAM t_b_359=3596.666667ns
.PARAM t_b_360=3609.98ns
.PARAM t_b_361=3616.666667ns
.PARAM t_b_362=3629.981ns
.PARAM t_b_363=3636.666667ns
.PARAM t_b_364=3649.982ns
.PARAM t_b_365=3656.666667ns
.PARAM t_b_366=3669.983ns
.PARAM t_b_367=3676.666667ns
.PARAM t_b_368=3689.984ns
.PARAM t_b_369=3696.666667ns
.PARAM t_b_370=3709.985ns
.PARAM t_b_371=3716.666667ns
.PARAM t_b_372=3729.986ns
.PARAM t_b_373=3736.666667ns
.PARAM t_b_374=3749.987ns
.PARAM t_b_375=3756.666667ns
.PARAM t_b_376=3769.988ns
.PARAM t_b_377=3776.666667ns
.PARAM t_b_378=3789.989ns
.PARAM t_b_379=3796.666667ns
.PARAM t_b_380=3809.99ns
.PARAM t_b_381=3816.666667ns
.PARAM t_b_382=3829.991ns
.PARAM t_b_383=3836.666667ns
.PARAM t_b_384=3849.992ns
.PARAM t_b_385=3856.666667ns
.PARAM t_b_386=3869.993ns
.PARAM t_b_387=3876.666667ns
.PARAM t_b_388=3889.994ns
.PARAM t_b_389=3896.666667ns
.PARAM t_b_390=3909.995ns
.PARAM t_b_391=3916.666667ns
.PARAM t_b_392=3929.996ns
.PARAM t_b_393=3936.666667ns
.PARAM t_b_394=3949.997ns
.PARAM t_b_395=3956.666667ns
.PARAM t_b_396=3969.998ns
.PARAM t_b_397=3976.666667ns
.PARAM t_b_398=3989.999ns
.PARAM t_b_399=3996.666667ns
.PARAM t_b_400=4010.0ns
.PARAM t_b_401=4016.666667ns
.PARAM t_b_402=4030.001ns
.PARAM t_b_403=4036.666667ns
.PARAM t_b_404=4050.002ns
.PARAM t_b_405=4056.666667ns
.PARAM t_b_406=4070.003ns
.PARAM t_b_407=4076.666667ns
.PARAM t_b_408=4090.004ns
.PARAM t_b_409=4096.666667ns
.PARAM t_b_410=4110.005ns
.PARAM t_b_411=4116.666667ns
.PARAM t_b_412=4130.006ns
.PARAM t_b_413=4136.666667ns
.PARAM t_b_414=4150.007ns
.PARAM t_b_415=4156.666667ns
.PARAM t_b_416=4170.008ns
.PARAM t_b_417=4176.666667ns
.PARAM t_b_418=4190.009ns
.PARAM t_b_419=4196.666667ns
.PARAM t_b_420=4210.01ns
.PARAM t_b_421=4216.666667ns
.PARAM t_b_422=4230.011ns
.PARAM t_b_423=4236.666667ns
.PARAM t_b_424=4250.012ns
.PARAM t_b_425=4256.666667ns
.PARAM t_b_426=4270.013ns
.PARAM t_b_427=4276.666667ns
.PARAM t_b_428=4290.014ns
.PARAM t_b_429=4296.666667ns
.PARAM t_b_430=4310.015ns
.PARAM t_b_431=4316.666667ns
.PARAM t_b_432=4330.016ns
.PARAM t_b_433=4336.666667ns
.PARAM t_b_434=4350.017ns
.PARAM t_b_435=4356.666667ns
.PARAM t_b_436=4370.018ns
.PARAM t_b_437=4376.666667ns
.PARAM t_b_438=4390.019ns
.PARAM t_b_439=4396.666667ns
.PARAM t_b_440=4410.02ns
.PARAM t_b_441=4416.666667ns
.PARAM t_b_442=4430.021ns
.PARAM t_b_443=4436.666667ns
.PARAM t_b_444=4450.022ns
.PARAM t_b_445=4456.666667ns
.PARAM t_b_446=4470.023ns
.PARAM t_b_447=4476.666667ns
.PARAM t_b_448=4490.024ns
.PARAM t_b_449=4496.666667ns
.PARAM t_b_450=4510.025ns
.PARAM t_b_451=4516.666667ns
.PARAM t_b_452=4530.026ns
.PARAM t_b_453=4536.666667ns
.PARAM t_b_454=4550.027ns
.PARAM t_b_455=4556.666667ns
.PARAM t_b_456=4570.028ns
.PARAM t_b_457=4576.666667ns
.PARAM t_b_458=4590.029ns
.PARAM t_b_459=4596.666667ns
.PARAM t_b_460=4610.03ns
.PARAM t_b_461=4616.666667ns
.PARAM t_b_462=4630.031ns
.PARAM t_b_463=4636.666667ns
.PARAM t_b_464=4650.032ns
.PARAM t_b_465=4656.666667ns
.PARAM t_b_466=4670.033ns
.PARAM t_b_467=4676.666667ns
.PARAM t_b_468=4690.034ns
.PARAM t_b_469=4696.666667ns
.PARAM t_b_470=4710.035ns
.PARAM t_b_471=4716.666667ns
.PARAM t_b_472=4730.036ns
.PARAM t_b_473=4736.666667ns
.PARAM t_b_474=4750.037ns
.PARAM t_b_475=4756.666667ns
.PARAM t_b_476=4770.038ns
.PARAM t_b_477=4776.666667ns
.PARAM t_b_478=4790.039ns
.PARAM t_b_479=4796.666667ns
.PARAM t_b_480=4810.04ns
.PARAM t_b_481=4816.666667ns
.PARAM t_b_482=4830.041ns
.PARAM t_b_483=4836.666667ns
.PARAM t_b_484=4850.042ns
.PARAM t_b_485=4856.666667ns
.PARAM t_b_486=4870.043ns
.PARAM t_b_487=4876.666667ns
.PARAM t_b_488=4890.044ns
.PARAM t_b_489=4896.666667ns
.PARAM t_b_490=4910.045ns
.PARAM t_b_491=4916.666667ns
.PARAM t_b_492=4930.046ns
.PARAM t_b_493=4936.666667ns
.PARAM t_b_494=4950.047ns
.PARAM t_b_495=4956.666667ns
.PARAM t_b_496=4970.048ns
.PARAM t_b_497=4976.666667ns
.PARAM t_b_498=4990.049ns
.PARAM t_b_499=4996.666667ns
.PARAM t_b_500=5010.05ns
.PARAM t_b_501=5016.666667ns
.PARAM t_b_502=5030.051ns
.PARAM t_b_503=5036.666667ns
.PARAM t_b_504=5050.052ns
.PARAM t_b_505=5056.666667ns
.PARAM t_b_506=5070.053ns
.PARAM t_b_507=5076.666667ns
.PARAM t_b_508=5090.054ns
.PARAM t_b_509=5096.666667ns
.PARAM t_b_510=5110.055ns
.PARAM t_b_511=5116.666667ns
.PARAM t_b_512=5130.056ns
.PARAM t_b_513=5136.666667ns
.PARAM t_b_514=5150.057ns
.PARAM t_b_515=5156.666667ns
.PARAM t_b_516=5170.058ns
.PARAM t_b_517=5176.666667ns
.PARAM t_b_518=5190.059ns
.PARAM t_b_519=5196.666667ns
.PARAM t_b_520=5210.06ns
.PARAM t_b_521=5216.666667ns
.PARAM t_b_522=5230.061ns
.PARAM t_b_523=5236.666667ns
.PARAM t_b_524=5250.062ns
.PARAM t_b_525=5256.666667ns
.PARAM t_b_526=5270.063ns
.PARAM t_b_527=5276.666667ns
.PARAM t_b_528=5290.064ns
.PARAM t_b_529=5296.666667ns
.PARAM t_b_530=5310.065ns
.PARAM t_b_531=5316.666667ns
.PARAM t_b_532=5330.066ns
.PARAM t_b_533=5336.666667ns
.PARAM t_b_534=5350.067ns
.PARAM t_b_535=5356.666667ns
.PARAM t_b_536=5370.068ns
.PARAM t_b_537=5376.666667ns
.PARAM t_b_538=5390.069ns
.PARAM t_b_539=5396.666667ns
.PARAM t_b_540=5410.07ns
.PARAM t_b_541=5416.666667ns
.PARAM t_b_542=5430.071ns
.PARAM t_b_543=5436.666667ns
.PARAM t_b_544=5450.072ns
.PARAM t_b_545=5456.666667ns
.PARAM t_b_546=5470.073ns
.PARAM t_b_547=5476.666667ns
.PARAM t_b_548=5490.074ns
.PARAM t_b_549=5496.666667ns
.PARAM t_b_550=5510.075ns
.PARAM t_b_551=5516.666667ns
.PARAM t_b_552=5530.076ns
.PARAM t_b_553=5536.666667ns
.PARAM t_b_554=5550.077ns
.PARAM t_b_555=5556.666667ns
.PARAM t_b_556=5570.078ns
.PARAM t_b_557=5576.666667ns
.PARAM t_b_558=5590.079ns
.PARAM t_b_559=5596.666667ns
.PARAM t_b_560=5610.08ns
.PARAM t_b_561=5616.666667ns
.PARAM t_b_562=5630.081ns
.PARAM t_b_563=5636.666667ns
.PARAM t_b_564=5650.082ns
.PARAM t_b_565=5656.666667ns
.PARAM t_b_566=5670.083ns
.PARAM t_b_567=5676.666667ns
.PARAM t_b_568=5690.084ns
.PARAM t_b_569=5696.666667ns
.PARAM t_b_570=5710.085ns
.PARAM t_b_571=5716.666667ns
.PARAM t_b_572=5730.086ns
.PARAM t_b_573=5736.666667ns
.PARAM t_b_574=5750.087ns
.PARAM t_b_575=5756.666667ns
.PARAM t_b_576=5770.088ns
.PARAM t_b_577=5776.666667ns
.PARAM t_b_578=5790.089ns
.PARAM t_b_579=5796.666667ns
.PARAM t_b_580=5810.09ns
.PARAM t_b_581=5816.666667ns
.PARAM t_b_582=5830.091ns
.PARAM t_b_583=5836.666667ns
.PARAM t_b_584=5850.092ns
.PARAM t_b_585=5856.666667ns
.PARAM t_b_586=5870.093ns
.PARAM t_b_587=5876.666667ns
.PARAM t_b_588=5890.094ns
.PARAM t_b_589=5896.666667ns
.PARAM t_b_590=5910.095ns
.PARAM t_b_591=5916.666667ns
.PARAM t_b_592=5930.096ns
.PARAM t_b_593=5936.666667ns
.PARAM t_b_594=5950.097ns
.PARAM t_b_595=5956.666667ns
.PARAM t_b_596=5970.098ns
.PARAM t_b_597=5976.666667ns
.PARAM t_b_598=5990.099ns
.PARAM t_b_599=5996.666667ns
.PARAM t_b_600=6010.1ns
.PARAM t_b_601=6016.666667ns
.PARAM t_b_602=6030.101ns
.PARAM t_b_603=6036.666667ns
.PARAM t_b_604=6050.102ns
.PARAM t_b_605=6056.666667ns
.PARAM t_b_606=6070.103ns
.PARAM t_b_607=6076.666667ns
.PARAM t_b_608=6090.104ns
.PARAM t_b_609=6096.666667ns
.PARAM t_b_610=6110.105ns
.PARAM t_b_611=6116.666667ns
.PARAM t_b_612=6130.106ns
.PARAM t_b_613=6136.666667ns
.PARAM t_b_614=6150.107ns
.PARAM t_b_615=6156.666667ns
.PARAM t_b_616=6170.108ns
.PARAM t_b_617=6176.666667ns
.PARAM t_b_618=6190.109ns
.PARAM t_b_619=6196.666667ns
.PARAM t_b_620=6210.11ns
.PARAM t_b_621=6216.666667ns
.PARAM t_b_622=6230.111ns
.PARAM t_b_623=6236.666667ns
.PARAM t_b_624=6250.112ns
.PARAM t_b_625=6256.666667ns
.PARAM t_b_626=6270.113ns
.PARAM t_b_627=6276.666667ns
.PARAM t_b_628=6290.114ns
.PARAM t_b_629=6296.666667ns
.PARAM t_b_630=6310.115ns
.PARAM t_b_631=6316.666667ns
.PARAM t_b_632=6330.116ns
.PARAM t_b_633=6336.666667ns
.PARAM t_b_634=6350.117ns
.PARAM t_b_635=6356.666667ns
.PARAM t_b_636=6370.118ns
.PARAM t_b_637=6376.666667ns
.PARAM t_b_638=6390.119ns
.PARAM t_b_639=6396.666667ns
.PARAM t_b_640=6410.12ns
.PARAM t_b_641=6416.666667ns
.PARAM t_b_642=6430.121ns
.PARAM t_b_643=6436.666667ns
.PARAM t_b_644=6450.122ns
.PARAM t_b_645=6456.666667ns
.PARAM t_b_646=6470.123ns
.PARAM t_b_647=6476.666667ns
.PARAM t_b_648=6490.124ns
.PARAM t_b_649=6496.666667ns
.PARAM t_b_650=6510.125ns
.PARAM t_b_651=6516.666667ns
.PARAM t_b_652=6530.126ns
.PARAM t_b_653=6536.666667ns
.PARAM t_b_654=6550.127ns
.PARAM t_b_655=6556.666667ns
.PARAM t_b_656=6570.128ns
.PARAM t_b_657=6576.666667ns
.PARAM t_b_658=6590.129ns
.PARAM t_b_659=6596.666667ns
.PARAM t_b_660=6610.13ns
.PARAM t_b_661=6616.666667ns
.PARAM t_b_662=6630.131ns
.PARAM t_b_663=6636.666667ns
.PARAM t_b_664=6650.132ns
.PARAM t_b_665=6656.666667ns
.PARAM t_b_666=6670.133ns
.PARAM t_b_667=6676.666667ns
.PARAM t_b_668=6690.134ns
.PARAM t_b_669=6696.666667ns
.PARAM t_b_670=6710.135ns
.PARAM t_b_671=6716.666667ns
.PARAM t_b_672=6730.136ns
.PARAM t_b_673=6736.666667ns
.PARAM t_b_674=6750.137ns
.PARAM t_b_675=6756.666667ns
.PARAM t_b_676=6770.138ns
.PARAM t_b_677=6776.666667ns
.PARAM t_b_678=6790.139ns
.PARAM t_b_679=6796.666667ns
.PARAM t_b_680=6810.14ns
.PARAM t_b_681=6816.666667ns
.PARAM t_b_682=6830.141ns
.PARAM t_b_683=6836.666667ns
.PARAM t_b_684=6850.142ns
.PARAM t_b_685=6856.666667ns
.PARAM t_b_686=6870.143ns
.PARAM t_b_687=6876.666667ns
.PARAM t_b_688=6890.144ns
.PARAM t_b_689=6896.666667ns
.PARAM t_b_690=6910.145ns
.PARAM t_b_691=6916.666667ns
.PARAM t_b_692=6930.146ns
.PARAM t_b_693=6936.666667ns
.PARAM t_b_694=6950.147ns
.PARAM t_b_695=6956.666667ns
.PARAM t_b_696=6970.148ns
.PARAM t_b_697=6976.666667ns
.PARAM t_b_698=6990.149ns
.PARAM t_b_699=6996.666667ns
.PARAM t_b_700=7010.15ns
.PARAM t_b_701=7016.666667ns
.PARAM t_b_702=7030.151ns
.PARAM t_b_703=7036.666667ns
.PARAM t_b_704=7050.152ns
.PARAM t_b_705=7056.666667ns
.PARAM t_b_706=7070.153ns
.PARAM t_b_707=7076.666667ns
.PARAM t_b_708=7090.154ns
.PARAM t_b_709=7096.666667ns
.PARAM t_b_710=7110.155ns
.PARAM t_b_711=7116.666667ns
.PARAM t_b_712=7130.156ns
.PARAM t_b_713=7136.666667ns
.PARAM t_b_714=7150.157ns
.PARAM t_b_715=7156.666667ns
.PARAM t_b_716=7170.158ns
.PARAM t_b_717=7176.666667ns
.PARAM t_b_718=7190.159ns
.PARAM t_b_719=7196.666667ns
.PARAM t_b_720=7210.16ns
.PARAM t_b_721=7216.666667ns
.PARAM t_b_722=7230.161ns
.PARAM t_b_723=7236.666667ns
.PARAM t_b_724=7250.162ns
.PARAM t_b_725=7256.666667ns
.PARAM t_b_726=7270.163ns
.PARAM t_b_727=7276.666667ns
.PARAM t_b_728=7290.164ns
.PARAM t_b_729=7296.666667ns
.PARAM t_b_730=7310.165ns
.PARAM t_b_731=7316.666667ns
.PARAM t_b_732=7330.166ns
.PARAM t_b_733=7336.666667ns
.PARAM t_b_734=7350.167ns
.PARAM t_b_735=7356.666667ns
.PARAM t_b_736=7370.168ns
.PARAM t_b_737=7376.666667ns
.PARAM t_b_738=7390.169ns
.PARAM t_b_739=7396.666667ns
.PARAM t_b_740=7410.17ns
.PARAM t_b_741=7416.666667ns
.PARAM t_b_742=7430.171ns
.PARAM t_b_743=7436.666667ns
.PARAM t_b_744=7450.172ns
.PARAM t_b_745=7456.666667ns
.PARAM t_b_746=7470.173ns
.PARAM t_b_747=7476.666667ns
.PARAM t_b_748=7490.174ns
.PARAM t_b_749=7496.666667ns
.PARAM t_b_750=7510.175ns
.PARAM t_b_751=7516.666667ns
.PARAM t_b_752=7530.176ns
.PARAM t_b_753=7536.666667ns
.PARAM t_b_754=7550.177ns
.PARAM t_b_755=7556.666667ns
.PARAM t_b_756=7570.178ns
.PARAM t_b_757=7576.666667ns
.PARAM t_b_758=7590.179ns
.PARAM t_b_759=7596.666667ns
.PARAM t_b_760=7610.18ns
.PARAM t_b_761=7616.666667ns
.PARAM t_b_762=7630.181ns
.PARAM t_b_763=7636.666667ns
.PARAM t_b_764=7650.182ns
.PARAM t_b_765=7656.666667ns
.PARAM t_b_766=7670.183ns
.PARAM t_b_767=7676.666667ns
.PARAM t_b_768=7690.184ns
.PARAM t_b_769=7696.666667ns
.PARAM t_b_770=7710.185ns
.PARAM t_b_771=7716.666667ns
.PARAM t_b_772=7730.186ns
.PARAM t_b_773=7736.666667ns
.PARAM t_b_774=7750.187ns
.PARAM t_b_775=7756.666667ns
.PARAM t_b_776=7770.188ns
.PARAM t_b_777=7776.666667ns
.PARAM t_b_778=7790.189ns
.PARAM t_b_779=7796.666667ns
.PARAM t_b_780=7810.19ns
.PARAM t_b_781=7816.666667ns
.PARAM t_b_782=7830.191ns
.PARAM t_b_783=7836.666667ns
.PARAM t_b_784=7850.192ns
.PARAM t_b_785=7856.666667ns
.PARAM t_b_786=7870.193ns
.PARAM t_b_787=7876.666667ns
.PARAM t_b_788=7890.194ns
.PARAM t_b_789=7896.666667ns
.PARAM t_b_790=7910.195ns
.PARAM t_b_791=7916.666667ns
.PARAM t_b_792=7930.196ns
.PARAM t_b_793=7936.666667ns
.PARAM t_b_794=7950.197ns
.PARAM t_b_795=7956.666667ns
.PARAM t_b_796=7970.198ns
.PARAM t_b_797=7976.666667ns
.PARAM t_b_798=7990.199ns
.PARAM t_b_799=7996.666667ns



VINA Input_A GND PWL 0ns baseVal t_init0 baseVal 't_init0+slope' peakVal t_init1 peakVal 't_init1+slope' baseVal
+ t_a_0 baseVal 't_a_0+slope' peakVal
+ t_a_1 peakVal 't_a_1+slope' baseVal
+ t_a_2 baseVal 't_a_2+slope' peakVal
+ t_a_3 peakVal 't_a_3+slope' baseVal
+ t_a_4 baseVal 't_a_4+slope' peakVal
+ t_a_5 peakVal 't_a_5+slope' baseVal
+ t_a_6 baseVal 't_a_6+slope' peakVal
+ t_a_7 peakVal 't_a_7+slope' baseVal
+ t_a_8 baseVal 't_a_8+slope' peakVal
+ t_a_9 peakVal 't_a_9+slope' baseVal
+ t_a_10 baseVal 't_a_10+slope' peakVal
+ t_a_11 peakVal 't_a_11+slope' baseVal
+ t_a_12 baseVal 't_a_12+slope' peakVal
+ t_a_13 peakVal 't_a_13+slope' baseVal
+ t_a_14 baseVal 't_a_14+slope' peakVal
+ t_a_15 peakVal 't_a_15+slope' baseVal
+ t_a_16 baseVal 't_a_16+slope' peakVal
+ t_a_17 peakVal 't_a_17+slope' baseVal
+ t_a_18 baseVal 't_a_18+slope' peakVal
+ t_a_19 peakVal 't_a_19+slope' baseVal
+ t_a_20 baseVal 't_a_20+slope' peakVal
+ t_a_21 peakVal 't_a_21+slope' baseVal
+ t_a_22 baseVal 't_a_22+slope' peakVal
+ t_a_23 peakVal 't_a_23+slope' baseVal
+ t_a_24 baseVal 't_a_24+slope' peakVal
+ t_a_25 peakVal 't_a_25+slope' baseVal
+ t_a_26 baseVal 't_a_26+slope' peakVal
+ t_a_27 peakVal 't_a_27+slope' baseVal
+ t_a_28 baseVal 't_a_28+slope' peakVal
+ t_a_29 peakVal 't_a_29+slope' baseVal
+ t_a_30 baseVal 't_a_30+slope' peakVal
+ t_a_31 peakVal 't_a_31+slope' baseVal
+ t_a_32 baseVal 't_a_32+slope' peakVal
+ t_a_33 peakVal 't_a_33+slope' baseVal
+ t_a_34 baseVal 't_a_34+slope' peakVal
+ t_a_35 peakVal 't_a_35+slope' baseVal
+ t_a_36 baseVal 't_a_36+slope' peakVal
+ t_a_37 peakVal 't_a_37+slope' baseVal
+ t_a_38 baseVal 't_a_38+slope' peakVal
+ t_a_39 peakVal 't_a_39+slope' baseVal
+ t_a_40 baseVal 't_a_40+slope' peakVal
+ t_a_41 peakVal 't_a_41+slope' baseVal
+ t_a_42 baseVal 't_a_42+slope' peakVal
+ t_a_43 peakVal 't_a_43+slope' baseVal
+ t_a_44 baseVal 't_a_44+slope' peakVal
+ t_a_45 peakVal 't_a_45+slope' baseVal
+ t_a_46 baseVal 't_a_46+slope' peakVal
+ t_a_47 peakVal 't_a_47+slope' baseVal
+ t_a_48 baseVal 't_a_48+slope' peakVal
+ t_a_49 peakVal 't_a_49+slope' baseVal
+ t_a_50 baseVal 't_a_50+slope' peakVal
+ t_a_51 peakVal 't_a_51+slope' baseVal
+ t_a_52 baseVal 't_a_52+slope' peakVal
+ t_a_53 peakVal 't_a_53+slope' baseVal
+ t_a_54 baseVal 't_a_54+slope' peakVal
+ t_a_55 peakVal 't_a_55+slope' baseVal
+ t_a_56 baseVal 't_a_56+slope' peakVal
+ t_a_57 peakVal 't_a_57+slope' baseVal
+ t_a_58 baseVal 't_a_58+slope' peakVal
+ t_a_59 peakVal 't_a_59+slope' baseVal
+ t_a_60 baseVal 't_a_60+slope' peakVal
+ t_a_61 peakVal 't_a_61+slope' baseVal
+ t_a_62 baseVal 't_a_62+slope' peakVal
+ t_a_63 peakVal 't_a_63+slope' baseVal
+ t_a_64 baseVal 't_a_64+slope' peakVal
+ t_a_65 peakVal 't_a_65+slope' baseVal
+ t_a_66 baseVal 't_a_66+slope' peakVal
+ t_a_67 peakVal 't_a_67+slope' baseVal
+ t_a_68 baseVal 't_a_68+slope' peakVal
+ t_a_69 peakVal 't_a_69+slope' baseVal
+ t_a_70 baseVal 't_a_70+slope' peakVal
+ t_a_71 peakVal 't_a_71+slope' baseVal
+ t_a_72 baseVal 't_a_72+slope' peakVal
+ t_a_73 peakVal 't_a_73+slope' baseVal
+ t_a_74 baseVal 't_a_74+slope' peakVal
+ t_a_75 peakVal 't_a_75+slope' baseVal
+ t_a_76 baseVal 't_a_76+slope' peakVal
+ t_a_77 peakVal 't_a_77+slope' baseVal
+ t_a_78 baseVal 't_a_78+slope' peakVal
+ t_a_79 peakVal 't_a_79+slope' baseVal
+ t_a_80 baseVal 't_a_80+slope' peakVal
+ t_a_81 peakVal 't_a_81+slope' baseVal
+ t_a_82 baseVal 't_a_82+slope' peakVal
+ t_a_83 peakVal 't_a_83+slope' baseVal
+ t_a_84 baseVal 't_a_84+slope' peakVal
+ t_a_85 peakVal 't_a_85+slope' baseVal
+ t_a_86 baseVal 't_a_86+slope' peakVal
+ t_a_87 peakVal 't_a_87+slope' baseVal
+ t_a_88 baseVal 't_a_88+slope' peakVal
+ t_a_89 peakVal 't_a_89+slope' baseVal
+ t_a_90 baseVal 't_a_90+slope' peakVal
+ t_a_91 peakVal 't_a_91+slope' baseVal
+ t_a_92 baseVal 't_a_92+slope' peakVal
+ t_a_93 peakVal 't_a_93+slope' baseVal
+ t_a_94 baseVal 't_a_94+slope' peakVal
+ t_a_95 peakVal 't_a_95+slope' baseVal
+ t_a_96 baseVal 't_a_96+slope' peakVal
+ t_a_97 peakVal 't_a_97+slope' baseVal
+ t_a_98 baseVal 't_a_98+slope' peakVal
+ t_a_99 peakVal 't_a_99+slope' baseVal
+ t_a_100 baseVal 't_a_100+slope' peakVal
+ t_a_101 peakVal 't_a_101+slope' baseVal
+ t_a_102 baseVal 't_a_102+slope' peakVal
+ t_a_103 peakVal 't_a_103+slope' baseVal
+ t_a_104 baseVal 't_a_104+slope' peakVal
+ t_a_105 peakVal 't_a_105+slope' baseVal
+ t_a_106 baseVal 't_a_106+slope' peakVal
+ t_a_107 peakVal 't_a_107+slope' baseVal
+ t_a_108 baseVal 't_a_108+slope' peakVal
+ t_a_109 peakVal 't_a_109+slope' baseVal
+ t_a_110 baseVal 't_a_110+slope' peakVal
+ t_a_111 peakVal 't_a_111+slope' baseVal
+ t_a_112 baseVal 't_a_112+slope' peakVal
+ t_a_113 peakVal 't_a_113+slope' baseVal
+ t_a_114 baseVal 't_a_114+slope' peakVal
+ t_a_115 peakVal 't_a_115+slope' baseVal
+ t_a_116 baseVal 't_a_116+slope' peakVal
+ t_a_117 peakVal 't_a_117+slope' baseVal
+ t_a_118 baseVal 't_a_118+slope' peakVal
+ t_a_119 peakVal 't_a_119+slope' baseVal
+ t_a_120 baseVal 't_a_120+slope' peakVal
+ t_a_121 peakVal 't_a_121+slope' baseVal
+ t_a_122 baseVal 't_a_122+slope' peakVal
+ t_a_123 peakVal 't_a_123+slope' baseVal
+ t_a_124 baseVal 't_a_124+slope' peakVal
+ t_a_125 peakVal 't_a_125+slope' baseVal
+ t_a_126 baseVal 't_a_126+slope' peakVal
+ t_a_127 peakVal 't_a_127+slope' baseVal
+ t_a_128 baseVal 't_a_128+slope' peakVal
+ t_a_129 peakVal 't_a_129+slope' baseVal
+ t_a_130 baseVal 't_a_130+slope' peakVal
+ t_a_131 peakVal 't_a_131+slope' baseVal
+ t_a_132 baseVal 't_a_132+slope' peakVal
+ t_a_133 peakVal 't_a_133+slope' baseVal
+ t_a_134 baseVal 't_a_134+slope' peakVal
+ t_a_135 peakVal 't_a_135+slope' baseVal
+ t_a_136 baseVal 't_a_136+slope' peakVal
+ t_a_137 peakVal 't_a_137+slope' baseVal
+ t_a_138 baseVal 't_a_138+slope' peakVal
+ t_a_139 peakVal 't_a_139+slope' baseVal
+ t_a_140 baseVal 't_a_140+slope' peakVal
+ t_a_141 peakVal 't_a_141+slope' baseVal
+ t_a_142 baseVal 't_a_142+slope' peakVal
+ t_a_143 peakVal 't_a_143+slope' baseVal
+ t_a_144 baseVal 't_a_144+slope' peakVal
+ t_a_145 peakVal 't_a_145+slope' baseVal
+ t_a_146 baseVal 't_a_146+slope' peakVal
+ t_a_147 peakVal 't_a_147+slope' baseVal
+ t_a_148 baseVal 't_a_148+slope' peakVal
+ t_a_149 peakVal 't_a_149+slope' baseVal
+ t_a_150 baseVal 't_a_150+slope' peakVal
+ t_a_151 peakVal 't_a_151+slope' baseVal
+ t_a_152 baseVal 't_a_152+slope' peakVal
+ t_a_153 peakVal 't_a_153+slope' baseVal
+ t_a_154 baseVal 't_a_154+slope' peakVal
+ t_a_155 peakVal 't_a_155+slope' baseVal
+ t_a_156 baseVal 't_a_156+slope' peakVal
+ t_a_157 peakVal 't_a_157+slope' baseVal
+ t_a_158 baseVal 't_a_158+slope' peakVal
+ t_a_159 peakVal 't_a_159+slope' baseVal
+ t_a_160 baseVal 't_a_160+slope' peakVal
+ t_a_161 peakVal 't_a_161+slope' baseVal
+ t_a_162 baseVal 't_a_162+slope' peakVal
+ t_a_163 peakVal 't_a_163+slope' baseVal
+ t_a_164 baseVal 't_a_164+slope' peakVal
+ t_a_165 peakVal 't_a_165+slope' baseVal
+ t_a_166 baseVal 't_a_166+slope' peakVal
+ t_a_167 peakVal 't_a_167+slope' baseVal
+ t_a_168 baseVal 't_a_168+slope' peakVal
+ t_a_169 peakVal 't_a_169+slope' baseVal
+ t_a_170 baseVal 't_a_170+slope' peakVal
+ t_a_171 peakVal 't_a_171+slope' baseVal
+ t_a_172 baseVal 't_a_172+slope' peakVal
+ t_a_173 peakVal 't_a_173+slope' baseVal
+ t_a_174 baseVal 't_a_174+slope' peakVal
+ t_a_175 peakVal 't_a_175+slope' baseVal
+ t_a_176 baseVal 't_a_176+slope' peakVal
+ t_a_177 peakVal 't_a_177+slope' baseVal
+ t_a_178 baseVal 't_a_178+slope' peakVal
+ t_a_179 peakVal 't_a_179+slope' baseVal
+ t_a_180 baseVal 't_a_180+slope' peakVal
+ t_a_181 peakVal 't_a_181+slope' baseVal
+ t_a_182 baseVal 't_a_182+slope' peakVal
+ t_a_183 peakVal 't_a_183+slope' baseVal
+ t_a_184 baseVal 't_a_184+slope' peakVal
+ t_a_185 peakVal 't_a_185+slope' baseVal
+ t_a_186 baseVal 't_a_186+slope' peakVal
+ t_a_187 peakVal 't_a_187+slope' baseVal
+ t_a_188 baseVal 't_a_188+slope' peakVal
+ t_a_189 peakVal 't_a_189+slope' baseVal
+ t_a_190 baseVal 't_a_190+slope' peakVal
+ t_a_191 peakVal 't_a_191+slope' baseVal
+ t_a_192 baseVal 't_a_192+slope' peakVal
+ t_a_193 peakVal 't_a_193+slope' baseVal
+ t_a_194 baseVal 't_a_194+slope' peakVal
+ t_a_195 peakVal 't_a_195+slope' baseVal
+ t_a_196 baseVal 't_a_196+slope' peakVal
+ t_a_197 peakVal 't_a_197+slope' baseVal
+ t_a_198 baseVal 't_a_198+slope' peakVal
+ t_a_199 peakVal 't_a_199+slope' baseVal
+ t_a_200 baseVal 't_a_200+slope' peakVal
+ t_a_201 peakVal 't_a_201+slope' baseVal
+ t_a_202 baseVal 't_a_202+slope' peakVal
+ t_a_203 peakVal 't_a_203+slope' baseVal
+ t_a_204 baseVal 't_a_204+slope' peakVal
+ t_a_205 peakVal 't_a_205+slope' baseVal
+ t_a_206 baseVal 't_a_206+slope' peakVal
+ t_a_207 peakVal 't_a_207+slope' baseVal
+ t_a_208 baseVal 't_a_208+slope' peakVal
+ t_a_209 peakVal 't_a_209+slope' baseVal
+ t_a_210 baseVal 't_a_210+slope' peakVal
+ t_a_211 peakVal 't_a_211+slope' baseVal
+ t_a_212 baseVal 't_a_212+slope' peakVal
+ t_a_213 peakVal 't_a_213+slope' baseVal
+ t_a_214 baseVal 't_a_214+slope' peakVal
+ t_a_215 peakVal 't_a_215+slope' baseVal
+ t_a_216 baseVal 't_a_216+slope' peakVal
+ t_a_217 peakVal 't_a_217+slope' baseVal
+ t_a_218 baseVal 't_a_218+slope' peakVal
+ t_a_219 peakVal 't_a_219+slope' baseVal
+ t_a_220 baseVal 't_a_220+slope' peakVal
+ t_a_221 peakVal 't_a_221+slope' baseVal
+ t_a_222 baseVal 't_a_222+slope' peakVal
+ t_a_223 peakVal 't_a_223+slope' baseVal
+ t_a_224 baseVal 't_a_224+slope' peakVal
+ t_a_225 peakVal 't_a_225+slope' baseVal
+ t_a_226 baseVal 't_a_226+slope' peakVal
+ t_a_227 peakVal 't_a_227+slope' baseVal
+ t_a_228 baseVal 't_a_228+slope' peakVal
+ t_a_229 peakVal 't_a_229+slope' baseVal
+ t_a_230 baseVal 't_a_230+slope' peakVal
+ t_a_231 peakVal 't_a_231+slope' baseVal
+ t_a_232 baseVal 't_a_232+slope' peakVal
+ t_a_233 peakVal 't_a_233+slope' baseVal
+ t_a_234 baseVal 't_a_234+slope' peakVal
+ t_a_235 peakVal 't_a_235+slope' baseVal
+ t_a_236 baseVal 't_a_236+slope' peakVal
+ t_a_237 peakVal 't_a_237+slope' baseVal
+ t_a_238 baseVal 't_a_238+slope' peakVal
+ t_a_239 peakVal 't_a_239+slope' baseVal
+ t_a_240 baseVal 't_a_240+slope' peakVal
+ t_a_241 peakVal 't_a_241+slope' baseVal
+ t_a_242 baseVal 't_a_242+slope' peakVal
+ t_a_243 peakVal 't_a_243+slope' baseVal
+ t_a_244 baseVal 't_a_244+slope' peakVal
+ t_a_245 peakVal 't_a_245+slope' baseVal
+ t_a_246 baseVal 't_a_246+slope' peakVal
+ t_a_247 peakVal 't_a_247+slope' baseVal
+ t_a_248 baseVal 't_a_248+slope' peakVal
+ t_a_249 peakVal 't_a_249+slope' baseVal
+ t_a_250 baseVal 't_a_250+slope' peakVal
+ t_a_251 peakVal 't_a_251+slope' baseVal
+ t_a_252 baseVal 't_a_252+slope' peakVal
+ t_a_253 peakVal 't_a_253+slope' baseVal
+ t_a_254 baseVal 't_a_254+slope' peakVal
+ t_a_255 peakVal 't_a_255+slope' baseVal
+ t_a_256 baseVal 't_a_256+slope' peakVal
+ t_a_257 peakVal 't_a_257+slope' baseVal
+ t_a_258 baseVal 't_a_258+slope' peakVal
+ t_a_259 peakVal 't_a_259+slope' baseVal
+ t_a_260 baseVal 't_a_260+slope' peakVal
+ t_a_261 peakVal 't_a_261+slope' baseVal
+ t_a_262 baseVal 't_a_262+slope' peakVal
+ t_a_263 peakVal 't_a_263+slope' baseVal
+ t_a_264 baseVal 't_a_264+slope' peakVal
+ t_a_265 peakVal 't_a_265+slope' baseVal
+ t_a_266 baseVal 't_a_266+slope' peakVal
+ t_a_267 peakVal 't_a_267+slope' baseVal
+ t_a_268 baseVal 't_a_268+slope' peakVal
+ t_a_269 peakVal 't_a_269+slope' baseVal
+ t_a_270 baseVal 't_a_270+slope' peakVal
+ t_a_271 peakVal 't_a_271+slope' baseVal
+ t_a_272 baseVal 't_a_272+slope' peakVal
+ t_a_273 peakVal 't_a_273+slope' baseVal
+ t_a_274 baseVal 't_a_274+slope' peakVal
+ t_a_275 peakVal 't_a_275+slope' baseVal
+ t_a_276 baseVal 't_a_276+slope' peakVal
+ t_a_277 peakVal 't_a_277+slope' baseVal
+ t_a_278 baseVal 't_a_278+slope' peakVal
+ t_a_279 peakVal 't_a_279+slope' baseVal
+ t_a_280 baseVal 't_a_280+slope' peakVal
+ t_a_281 peakVal 't_a_281+slope' baseVal
+ t_a_282 baseVal 't_a_282+slope' peakVal
+ t_a_283 peakVal 't_a_283+slope' baseVal
+ t_a_284 baseVal 't_a_284+slope' peakVal
+ t_a_285 peakVal 't_a_285+slope' baseVal
+ t_a_286 baseVal 't_a_286+slope' peakVal
+ t_a_287 peakVal 't_a_287+slope' baseVal
+ t_a_288 baseVal 't_a_288+slope' peakVal
+ t_a_289 peakVal 't_a_289+slope' baseVal
+ t_a_290 baseVal 't_a_290+slope' peakVal
+ t_a_291 peakVal 't_a_291+slope' baseVal
+ t_a_292 baseVal 't_a_292+slope' peakVal
+ t_a_293 peakVal 't_a_293+slope' baseVal
+ t_a_294 baseVal 't_a_294+slope' peakVal
+ t_a_295 peakVal 't_a_295+slope' baseVal
+ t_a_296 baseVal 't_a_296+slope' peakVal
+ t_a_297 peakVal 't_a_297+slope' baseVal
+ t_a_298 baseVal 't_a_298+slope' peakVal
+ t_a_299 peakVal 't_a_299+slope' baseVal
+ t_a_300 baseVal 't_a_300+slope' peakVal
+ t_a_301 peakVal 't_a_301+slope' baseVal
+ t_a_302 baseVal 't_a_302+slope' peakVal
+ t_a_303 peakVal 't_a_303+slope' baseVal
+ t_a_304 baseVal 't_a_304+slope' peakVal
+ t_a_305 peakVal 't_a_305+slope' baseVal
+ t_a_306 baseVal 't_a_306+slope' peakVal
+ t_a_307 peakVal 't_a_307+slope' baseVal
+ t_a_308 baseVal 't_a_308+slope' peakVal
+ t_a_309 peakVal 't_a_309+slope' baseVal
+ t_a_310 baseVal 't_a_310+slope' peakVal
+ t_a_311 peakVal 't_a_311+slope' baseVal
+ t_a_312 baseVal 't_a_312+slope' peakVal
+ t_a_313 peakVal 't_a_313+slope' baseVal
+ t_a_314 baseVal 't_a_314+slope' peakVal
+ t_a_315 peakVal 't_a_315+slope' baseVal
+ t_a_316 baseVal 't_a_316+slope' peakVal
+ t_a_317 peakVal 't_a_317+slope' baseVal
+ t_a_318 baseVal 't_a_318+slope' peakVal
+ t_a_319 peakVal 't_a_319+slope' baseVal
+ t_a_320 baseVal 't_a_320+slope' peakVal
+ t_a_321 peakVal 't_a_321+slope' baseVal
+ t_a_322 baseVal 't_a_322+slope' peakVal
+ t_a_323 peakVal 't_a_323+slope' baseVal
+ t_a_324 baseVal 't_a_324+slope' peakVal
+ t_a_325 peakVal 't_a_325+slope' baseVal
+ t_a_326 baseVal 't_a_326+slope' peakVal
+ t_a_327 peakVal 't_a_327+slope' baseVal
+ t_a_328 baseVal 't_a_328+slope' peakVal
+ t_a_329 peakVal 't_a_329+slope' baseVal
+ t_a_330 baseVal 't_a_330+slope' peakVal
+ t_a_331 peakVal 't_a_331+slope' baseVal
+ t_a_332 baseVal 't_a_332+slope' peakVal
+ t_a_333 peakVal 't_a_333+slope' baseVal
+ t_a_334 baseVal 't_a_334+slope' peakVal
+ t_a_335 peakVal 't_a_335+slope' baseVal
+ t_a_336 baseVal 't_a_336+slope' peakVal
+ t_a_337 peakVal 't_a_337+slope' baseVal
+ t_a_338 baseVal 't_a_338+slope' peakVal
+ t_a_339 peakVal 't_a_339+slope' baseVal
+ t_a_340 baseVal 't_a_340+slope' peakVal
+ t_a_341 peakVal 't_a_341+slope' baseVal
+ t_a_342 baseVal 't_a_342+slope' peakVal
+ t_a_343 peakVal 't_a_343+slope' baseVal
+ t_a_344 baseVal 't_a_344+slope' peakVal
+ t_a_345 peakVal 't_a_345+slope' baseVal
+ t_a_346 baseVal 't_a_346+slope' peakVal
+ t_a_347 peakVal 't_a_347+slope' baseVal
+ t_a_348 baseVal 't_a_348+slope' peakVal
+ t_a_349 peakVal 't_a_349+slope' baseVal
+ t_a_350 baseVal 't_a_350+slope' peakVal
+ t_a_351 peakVal 't_a_351+slope' baseVal
+ t_a_352 baseVal 't_a_352+slope' peakVal
+ t_a_353 peakVal 't_a_353+slope' baseVal
+ t_a_354 baseVal 't_a_354+slope' peakVal
+ t_a_355 peakVal 't_a_355+slope' baseVal
+ t_a_356 baseVal 't_a_356+slope' peakVal
+ t_a_357 peakVal 't_a_357+slope' baseVal
+ t_a_358 baseVal 't_a_358+slope' peakVal
+ t_a_359 peakVal 't_a_359+slope' baseVal
+ t_a_360 baseVal 't_a_360+slope' peakVal
+ t_a_361 peakVal 't_a_361+slope' baseVal
+ t_a_362 baseVal 't_a_362+slope' peakVal
+ t_a_363 peakVal 't_a_363+slope' baseVal
+ t_a_364 baseVal 't_a_364+slope' peakVal
+ t_a_365 peakVal 't_a_365+slope' baseVal
+ t_a_366 baseVal 't_a_366+slope' peakVal
+ t_a_367 peakVal 't_a_367+slope' baseVal
+ t_a_368 baseVal 't_a_368+slope' peakVal
+ t_a_369 peakVal 't_a_369+slope' baseVal
+ t_a_370 baseVal 't_a_370+slope' peakVal
+ t_a_371 peakVal 't_a_371+slope' baseVal
+ t_a_372 baseVal 't_a_372+slope' peakVal
+ t_a_373 peakVal 't_a_373+slope' baseVal
+ t_a_374 baseVal 't_a_374+slope' peakVal
+ t_a_375 peakVal 't_a_375+slope' baseVal
+ t_a_376 baseVal 't_a_376+slope' peakVal
+ t_a_377 peakVal 't_a_377+slope' baseVal
+ t_a_378 baseVal 't_a_378+slope' peakVal
+ t_a_379 peakVal 't_a_379+slope' baseVal
+ t_a_380 baseVal 't_a_380+slope' peakVal
+ t_a_381 peakVal 't_a_381+slope' baseVal
+ t_a_382 baseVal 't_a_382+slope' peakVal
+ t_a_383 peakVal 't_a_383+slope' baseVal
+ t_a_384 baseVal 't_a_384+slope' peakVal
+ t_a_385 peakVal 't_a_385+slope' baseVal
+ t_a_386 baseVal 't_a_386+slope' peakVal
+ t_a_387 peakVal 't_a_387+slope' baseVal
+ t_a_388 baseVal 't_a_388+slope' peakVal
+ t_a_389 peakVal 't_a_389+slope' baseVal
+ t_a_390 baseVal 't_a_390+slope' peakVal
+ t_a_391 peakVal 't_a_391+slope' baseVal
+ t_a_392 baseVal 't_a_392+slope' peakVal
+ t_a_393 peakVal 't_a_393+slope' baseVal
+ t_a_394 baseVal 't_a_394+slope' peakVal
+ t_a_395 peakVal 't_a_395+slope' baseVal
+ t_a_396 baseVal 't_a_396+slope' peakVal
+ t_a_397 peakVal 't_a_397+slope' baseVal
+ t_a_398 baseVal 't_a_398+slope' peakVal
+ t_a_399 peakVal 't_a_399+slope' baseVal
+ t_a_400 baseVal 't_a_400+slope' peakVal
+ t_a_401 peakVal 't_a_401+slope' baseVal
+ t_a_402 baseVal 't_a_402+slope' peakVal
+ t_a_403 peakVal 't_a_403+slope' baseVal
+ t_a_404 baseVal 't_a_404+slope' peakVal
+ t_a_405 peakVal 't_a_405+slope' baseVal
+ t_a_406 baseVal 't_a_406+slope' peakVal
+ t_a_407 peakVal 't_a_407+slope' baseVal
+ t_a_408 baseVal 't_a_408+slope' peakVal
+ t_a_409 peakVal 't_a_409+slope' baseVal
+ t_a_410 baseVal 't_a_410+slope' peakVal
+ t_a_411 peakVal 't_a_411+slope' baseVal
+ t_a_412 baseVal 't_a_412+slope' peakVal
+ t_a_413 peakVal 't_a_413+slope' baseVal
+ t_a_414 baseVal 't_a_414+slope' peakVal
+ t_a_415 peakVal 't_a_415+slope' baseVal
+ t_a_416 baseVal 't_a_416+slope' peakVal
+ t_a_417 peakVal 't_a_417+slope' baseVal
+ t_a_418 baseVal 't_a_418+slope' peakVal
+ t_a_419 peakVal 't_a_419+slope' baseVal
+ t_a_420 baseVal 't_a_420+slope' peakVal
+ t_a_421 peakVal 't_a_421+slope' baseVal
+ t_a_422 baseVal 't_a_422+slope' peakVal
+ t_a_423 peakVal 't_a_423+slope' baseVal
+ t_a_424 baseVal 't_a_424+slope' peakVal
+ t_a_425 peakVal 't_a_425+slope' baseVal
+ t_a_426 baseVal 't_a_426+slope' peakVal
+ t_a_427 peakVal 't_a_427+slope' baseVal
+ t_a_428 baseVal 't_a_428+slope' peakVal
+ t_a_429 peakVal 't_a_429+slope' baseVal
+ t_a_430 baseVal 't_a_430+slope' peakVal
+ t_a_431 peakVal 't_a_431+slope' baseVal
+ t_a_432 baseVal 't_a_432+slope' peakVal
+ t_a_433 peakVal 't_a_433+slope' baseVal
+ t_a_434 baseVal 't_a_434+slope' peakVal
+ t_a_435 peakVal 't_a_435+slope' baseVal
+ t_a_436 baseVal 't_a_436+slope' peakVal
+ t_a_437 peakVal 't_a_437+slope' baseVal
+ t_a_438 baseVal 't_a_438+slope' peakVal
+ t_a_439 peakVal 't_a_439+slope' baseVal
+ t_a_440 baseVal 't_a_440+slope' peakVal
+ t_a_441 peakVal 't_a_441+slope' baseVal
+ t_a_442 baseVal 't_a_442+slope' peakVal
+ t_a_443 peakVal 't_a_443+slope' baseVal
+ t_a_444 baseVal 't_a_444+slope' peakVal
+ t_a_445 peakVal 't_a_445+slope' baseVal
+ t_a_446 baseVal 't_a_446+slope' peakVal
+ t_a_447 peakVal 't_a_447+slope' baseVal
+ t_a_448 baseVal 't_a_448+slope' peakVal
+ t_a_449 peakVal 't_a_449+slope' baseVal
+ t_a_450 baseVal 't_a_450+slope' peakVal
+ t_a_451 peakVal 't_a_451+slope' baseVal
+ t_a_452 baseVal 't_a_452+slope' peakVal
+ t_a_453 peakVal 't_a_453+slope' baseVal
+ t_a_454 baseVal 't_a_454+slope' peakVal
+ t_a_455 peakVal 't_a_455+slope' baseVal
+ t_a_456 baseVal 't_a_456+slope' peakVal
+ t_a_457 peakVal 't_a_457+slope' baseVal
+ t_a_458 baseVal 't_a_458+slope' peakVal
+ t_a_459 peakVal 't_a_459+slope' baseVal
+ t_a_460 baseVal 't_a_460+slope' peakVal
+ t_a_461 peakVal 't_a_461+slope' baseVal
+ t_a_462 baseVal 't_a_462+slope' peakVal
+ t_a_463 peakVal 't_a_463+slope' baseVal
+ t_a_464 baseVal 't_a_464+slope' peakVal
+ t_a_465 peakVal 't_a_465+slope' baseVal
+ t_a_466 baseVal 't_a_466+slope' peakVal
+ t_a_467 peakVal 't_a_467+slope' baseVal
+ t_a_468 baseVal 't_a_468+slope' peakVal
+ t_a_469 peakVal 't_a_469+slope' baseVal
+ t_a_470 baseVal 't_a_470+slope' peakVal
+ t_a_471 peakVal 't_a_471+slope' baseVal
+ t_a_472 baseVal 't_a_472+slope' peakVal
+ t_a_473 peakVal 't_a_473+slope' baseVal
+ t_a_474 baseVal 't_a_474+slope' peakVal
+ t_a_475 peakVal 't_a_475+slope' baseVal
+ t_a_476 baseVal 't_a_476+slope' peakVal
+ t_a_477 peakVal 't_a_477+slope' baseVal
+ t_a_478 baseVal 't_a_478+slope' peakVal
+ t_a_479 peakVal 't_a_479+slope' baseVal
+ t_a_480 baseVal 't_a_480+slope' peakVal
+ t_a_481 peakVal 't_a_481+slope' baseVal
+ t_a_482 baseVal 't_a_482+slope' peakVal
+ t_a_483 peakVal 't_a_483+slope' baseVal
+ t_a_484 baseVal 't_a_484+slope' peakVal
+ t_a_485 peakVal 't_a_485+slope' baseVal
+ t_a_486 baseVal 't_a_486+slope' peakVal
+ t_a_487 peakVal 't_a_487+slope' baseVal
+ t_a_488 baseVal 't_a_488+slope' peakVal
+ t_a_489 peakVal 't_a_489+slope' baseVal
+ t_a_490 baseVal 't_a_490+slope' peakVal
+ t_a_491 peakVal 't_a_491+slope' baseVal
+ t_a_492 baseVal 't_a_492+slope' peakVal
+ t_a_493 peakVal 't_a_493+slope' baseVal
+ t_a_494 baseVal 't_a_494+slope' peakVal
+ t_a_495 peakVal 't_a_495+slope' baseVal
+ t_a_496 baseVal 't_a_496+slope' peakVal
+ t_a_497 peakVal 't_a_497+slope' baseVal
+ t_a_498 baseVal 't_a_498+slope' peakVal
+ t_a_499 peakVal 't_a_499+slope' baseVal
+ t_a_500 baseVal 't_a_500+slope' peakVal
+ t_a_501 peakVal 't_a_501+slope' baseVal
+ t_a_502 baseVal 't_a_502+slope' peakVal
+ t_a_503 peakVal 't_a_503+slope' baseVal
+ t_a_504 baseVal 't_a_504+slope' peakVal
+ t_a_505 peakVal 't_a_505+slope' baseVal
+ t_a_506 baseVal 't_a_506+slope' peakVal
+ t_a_507 peakVal 't_a_507+slope' baseVal
+ t_a_508 baseVal 't_a_508+slope' peakVal
+ t_a_509 peakVal 't_a_509+slope' baseVal
+ t_a_510 baseVal 't_a_510+slope' peakVal
+ t_a_511 peakVal 't_a_511+slope' baseVal
+ t_a_512 baseVal 't_a_512+slope' peakVal
+ t_a_513 peakVal 't_a_513+slope' baseVal
+ t_a_514 baseVal 't_a_514+slope' peakVal
+ t_a_515 peakVal 't_a_515+slope' baseVal
+ t_a_516 baseVal 't_a_516+slope' peakVal
+ t_a_517 peakVal 't_a_517+slope' baseVal
+ t_a_518 baseVal 't_a_518+slope' peakVal
+ t_a_519 peakVal 't_a_519+slope' baseVal
+ t_a_520 baseVal 't_a_520+slope' peakVal
+ t_a_521 peakVal 't_a_521+slope' baseVal
+ t_a_522 baseVal 't_a_522+slope' peakVal
+ t_a_523 peakVal 't_a_523+slope' baseVal
+ t_a_524 baseVal 't_a_524+slope' peakVal
+ t_a_525 peakVal 't_a_525+slope' baseVal
+ t_a_526 baseVal 't_a_526+slope' peakVal
+ t_a_527 peakVal 't_a_527+slope' baseVal
+ t_a_528 baseVal 't_a_528+slope' peakVal
+ t_a_529 peakVal 't_a_529+slope' baseVal
+ t_a_530 baseVal 't_a_530+slope' peakVal
+ t_a_531 peakVal 't_a_531+slope' baseVal
+ t_a_532 baseVal 't_a_532+slope' peakVal
+ t_a_533 peakVal 't_a_533+slope' baseVal
+ t_a_534 baseVal 't_a_534+slope' peakVal
+ t_a_535 peakVal 't_a_535+slope' baseVal
+ t_a_536 baseVal 't_a_536+slope' peakVal
+ t_a_537 peakVal 't_a_537+slope' baseVal
+ t_a_538 baseVal 't_a_538+slope' peakVal
+ t_a_539 peakVal 't_a_539+slope' baseVal
+ t_a_540 baseVal 't_a_540+slope' peakVal
+ t_a_541 peakVal 't_a_541+slope' baseVal
+ t_a_542 baseVal 't_a_542+slope' peakVal
+ t_a_543 peakVal 't_a_543+slope' baseVal
+ t_a_544 baseVal 't_a_544+slope' peakVal
+ t_a_545 peakVal 't_a_545+slope' baseVal
+ t_a_546 baseVal 't_a_546+slope' peakVal
+ t_a_547 peakVal 't_a_547+slope' baseVal
+ t_a_548 baseVal 't_a_548+slope' peakVal
+ t_a_549 peakVal 't_a_549+slope' baseVal
+ t_a_550 baseVal 't_a_550+slope' peakVal
+ t_a_551 peakVal 't_a_551+slope' baseVal
+ t_a_552 baseVal 't_a_552+slope' peakVal
+ t_a_553 peakVal 't_a_553+slope' baseVal
+ t_a_554 baseVal 't_a_554+slope' peakVal
+ t_a_555 peakVal 't_a_555+slope' baseVal
+ t_a_556 baseVal 't_a_556+slope' peakVal
+ t_a_557 peakVal 't_a_557+slope' baseVal
+ t_a_558 baseVal 't_a_558+slope' peakVal
+ t_a_559 peakVal 't_a_559+slope' baseVal
+ t_a_560 baseVal 't_a_560+slope' peakVal
+ t_a_561 peakVal 't_a_561+slope' baseVal
+ t_a_562 baseVal 't_a_562+slope' peakVal
+ t_a_563 peakVal 't_a_563+slope' baseVal
+ t_a_564 baseVal 't_a_564+slope' peakVal
+ t_a_565 peakVal 't_a_565+slope' baseVal
+ t_a_566 baseVal 't_a_566+slope' peakVal
+ t_a_567 peakVal 't_a_567+slope' baseVal
+ t_a_568 baseVal 't_a_568+slope' peakVal
+ t_a_569 peakVal 't_a_569+slope' baseVal
+ t_a_570 baseVal 't_a_570+slope' peakVal
+ t_a_571 peakVal 't_a_571+slope' baseVal
+ t_a_572 baseVal 't_a_572+slope' peakVal
+ t_a_573 peakVal 't_a_573+slope' baseVal
+ t_a_574 baseVal 't_a_574+slope' peakVal
+ t_a_575 peakVal 't_a_575+slope' baseVal
+ t_a_576 baseVal 't_a_576+slope' peakVal
+ t_a_577 peakVal 't_a_577+slope' baseVal
+ t_a_578 baseVal 't_a_578+slope' peakVal
+ t_a_579 peakVal 't_a_579+slope' baseVal
+ t_a_580 baseVal 't_a_580+slope' peakVal
+ t_a_581 peakVal 't_a_581+slope' baseVal
+ t_a_582 baseVal 't_a_582+slope' peakVal
+ t_a_583 peakVal 't_a_583+slope' baseVal
+ t_a_584 baseVal 't_a_584+slope' peakVal
+ t_a_585 peakVal 't_a_585+slope' baseVal
+ t_a_586 baseVal 't_a_586+slope' peakVal
+ t_a_587 peakVal 't_a_587+slope' baseVal
+ t_a_588 baseVal 't_a_588+slope' peakVal
+ t_a_589 peakVal 't_a_589+slope' baseVal
+ t_a_590 baseVal 't_a_590+slope' peakVal
+ t_a_591 peakVal 't_a_591+slope' baseVal
+ t_a_592 baseVal 't_a_592+slope' peakVal
+ t_a_593 peakVal 't_a_593+slope' baseVal
+ t_a_594 baseVal 't_a_594+slope' peakVal
+ t_a_595 peakVal 't_a_595+slope' baseVal
+ t_a_596 baseVal 't_a_596+slope' peakVal
+ t_a_597 peakVal 't_a_597+slope' baseVal
+ t_a_598 baseVal 't_a_598+slope' peakVal
+ t_a_599 peakVal 't_a_599+slope' baseVal
+ t_a_600 baseVal 't_a_600+slope' peakVal
+ t_a_601 peakVal 't_a_601+slope' baseVal
+ t_a_602 baseVal 't_a_602+slope' peakVal
+ t_a_603 peakVal 't_a_603+slope' baseVal
+ t_a_604 baseVal 't_a_604+slope' peakVal
+ t_a_605 peakVal 't_a_605+slope' baseVal
+ t_a_606 baseVal 't_a_606+slope' peakVal
+ t_a_607 peakVal 't_a_607+slope' baseVal
+ t_a_608 baseVal 't_a_608+slope' peakVal
+ t_a_609 peakVal 't_a_609+slope' baseVal
+ t_a_610 baseVal 't_a_610+slope' peakVal
+ t_a_611 peakVal 't_a_611+slope' baseVal
+ t_a_612 baseVal 't_a_612+slope' peakVal
+ t_a_613 peakVal 't_a_613+slope' baseVal
+ t_a_614 baseVal 't_a_614+slope' peakVal
+ t_a_615 peakVal 't_a_615+slope' baseVal
+ t_a_616 baseVal 't_a_616+slope' peakVal
+ t_a_617 peakVal 't_a_617+slope' baseVal
+ t_a_618 baseVal 't_a_618+slope' peakVal
+ t_a_619 peakVal 't_a_619+slope' baseVal
+ t_a_620 baseVal 't_a_620+slope' peakVal
+ t_a_621 peakVal 't_a_621+slope' baseVal
+ t_a_622 baseVal 't_a_622+slope' peakVal
+ t_a_623 peakVal 't_a_623+slope' baseVal
+ t_a_624 baseVal 't_a_624+slope' peakVal
+ t_a_625 peakVal 't_a_625+slope' baseVal
+ t_a_626 baseVal 't_a_626+slope' peakVal
+ t_a_627 peakVal 't_a_627+slope' baseVal
+ t_a_628 baseVal 't_a_628+slope' peakVal
+ t_a_629 peakVal 't_a_629+slope' baseVal
+ t_a_630 baseVal 't_a_630+slope' peakVal
+ t_a_631 peakVal 't_a_631+slope' baseVal
+ t_a_632 baseVal 't_a_632+slope' peakVal
+ t_a_633 peakVal 't_a_633+slope' baseVal
+ t_a_634 baseVal 't_a_634+slope' peakVal
+ t_a_635 peakVal 't_a_635+slope' baseVal
+ t_a_636 baseVal 't_a_636+slope' peakVal
+ t_a_637 peakVal 't_a_637+slope' baseVal
+ t_a_638 baseVal 't_a_638+slope' peakVal
+ t_a_639 peakVal 't_a_639+slope' baseVal
+ t_a_640 baseVal 't_a_640+slope' peakVal
+ t_a_641 peakVal 't_a_641+slope' baseVal
+ t_a_642 baseVal 't_a_642+slope' peakVal
+ t_a_643 peakVal 't_a_643+slope' baseVal
+ t_a_644 baseVal 't_a_644+slope' peakVal
+ t_a_645 peakVal 't_a_645+slope' baseVal
+ t_a_646 baseVal 't_a_646+slope' peakVal
+ t_a_647 peakVal 't_a_647+slope' baseVal
+ t_a_648 baseVal 't_a_648+slope' peakVal
+ t_a_649 peakVal 't_a_649+slope' baseVal
+ t_a_650 baseVal 't_a_650+slope' peakVal
+ t_a_651 peakVal 't_a_651+slope' baseVal
+ t_a_652 baseVal 't_a_652+slope' peakVal
+ t_a_653 peakVal 't_a_653+slope' baseVal
+ t_a_654 baseVal 't_a_654+slope' peakVal
+ t_a_655 peakVal 't_a_655+slope' baseVal
+ t_a_656 baseVal 't_a_656+slope' peakVal
+ t_a_657 peakVal 't_a_657+slope' baseVal
+ t_a_658 baseVal 't_a_658+slope' peakVal
+ t_a_659 peakVal 't_a_659+slope' baseVal
+ t_a_660 baseVal 't_a_660+slope' peakVal
+ t_a_661 peakVal 't_a_661+slope' baseVal
+ t_a_662 baseVal 't_a_662+slope' peakVal
+ t_a_663 peakVal 't_a_663+slope' baseVal
+ t_a_664 baseVal 't_a_664+slope' peakVal
+ t_a_665 peakVal 't_a_665+slope' baseVal
+ t_a_666 baseVal 't_a_666+slope' peakVal
+ t_a_667 peakVal 't_a_667+slope' baseVal
+ t_a_668 baseVal 't_a_668+slope' peakVal
+ t_a_669 peakVal 't_a_669+slope' baseVal
+ t_a_670 baseVal 't_a_670+slope' peakVal
+ t_a_671 peakVal 't_a_671+slope' baseVal
+ t_a_672 baseVal 't_a_672+slope' peakVal
+ t_a_673 peakVal 't_a_673+slope' baseVal
+ t_a_674 baseVal 't_a_674+slope' peakVal
+ t_a_675 peakVal 't_a_675+slope' baseVal
+ t_a_676 baseVal 't_a_676+slope' peakVal
+ t_a_677 peakVal 't_a_677+slope' baseVal
+ t_a_678 baseVal 't_a_678+slope' peakVal
+ t_a_679 peakVal 't_a_679+slope' baseVal
+ t_a_680 baseVal 't_a_680+slope' peakVal
+ t_a_681 peakVal 't_a_681+slope' baseVal
+ t_a_682 baseVal 't_a_682+slope' peakVal
+ t_a_683 peakVal 't_a_683+slope' baseVal
+ t_a_684 baseVal 't_a_684+slope' peakVal
+ t_a_685 peakVal 't_a_685+slope' baseVal
+ t_a_686 baseVal 't_a_686+slope' peakVal
+ t_a_687 peakVal 't_a_687+slope' baseVal
+ t_a_688 baseVal 't_a_688+slope' peakVal
+ t_a_689 peakVal 't_a_689+slope' baseVal
+ t_a_690 baseVal 't_a_690+slope' peakVal
+ t_a_691 peakVal 't_a_691+slope' baseVal
+ t_a_692 baseVal 't_a_692+slope' peakVal
+ t_a_693 peakVal 't_a_693+slope' baseVal
+ t_a_694 baseVal 't_a_694+slope' peakVal
+ t_a_695 peakVal 't_a_695+slope' baseVal
+ t_a_696 baseVal 't_a_696+slope' peakVal
+ t_a_697 peakVal 't_a_697+slope' baseVal
+ t_a_698 baseVal 't_a_698+slope' peakVal
+ t_a_699 peakVal 't_a_699+slope' baseVal
+ t_a_700 baseVal 't_a_700+slope' peakVal
+ t_a_701 peakVal 't_a_701+slope' baseVal
+ t_a_702 baseVal 't_a_702+slope' peakVal
+ t_a_703 peakVal 't_a_703+slope' baseVal
+ t_a_704 baseVal 't_a_704+slope' peakVal
+ t_a_705 peakVal 't_a_705+slope' baseVal
+ t_a_706 baseVal 't_a_706+slope' peakVal
+ t_a_707 peakVal 't_a_707+slope' baseVal
+ t_a_708 baseVal 't_a_708+slope' peakVal
+ t_a_709 peakVal 't_a_709+slope' baseVal
+ t_a_710 baseVal 't_a_710+slope' peakVal
+ t_a_711 peakVal 't_a_711+slope' baseVal
+ t_a_712 baseVal 't_a_712+slope' peakVal
+ t_a_713 peakVal 't_a_713+slope' baseVal
+ t_a_714 baseVal 't_a_714+slope' peakVal
+ t_a_715 peakVal 't_a_715+slope' baseVal
+ t_a_716 baseVal 't_a_716+slope' peakVal
+ t_a_717 peakVal 't_a_717+slope' baseVal
+ t_a_718 baseVal 't_a_718+slope' peakVal
+ t_a_719 peakVal 't_a_719+slope' baseVal
+ t_a_720 baseVal 't_a_720+slope' peakVal
+ t_a_721 peakVal 't_a_721+slope' baseVal
+ t_a_722 baseVal 't_a_722+slope' peakVal
+ t_a_723 peakVal 't_a_723+slope' baseVal
+ t_a_724 baseVal 't_a_724+slope' peakVal
+ t_a_725 peakVal 't_a_725+slope' baseVal
+ t_a_726 baseVal 't_a_726+slope' peakVal
+ t_a_727 peakVal 't_a_727+slope' baseVal
+ t_a_728 baseVal 't_a_728+slope' peakVal
+ t_a_729 peakVal 't_a_729+slope' baseVal
+ t_a_730 baseVal 't_a_730+slope' peakVal
+ t_a_731 peakVal 't_a_731+slope' baseVal
+ t_a_732 baseVal 't_a_732+slope' peakVal
+ t_a_733 peakVal 't_a_733+slope' baseVal
+ t_a_734 baseVal 't_a_734+slope' peakVal
+ t_a_735 peakVal 't_a_735+slope' baseVal
+ t_a_736 baseVal 't_a_736+slope' peakVal
+ t_a_737 peakVal 't_a_737+slope' baseVal
+ t_a_738 baseVal 't_a_738+slope' peakVal
+ t_a_739 peakVal 't_a_739+slope' baseVal
+ t_a_740 baseVal 't_a_740+slope' peakVal
+ t_a_741 peakVal 't_a_741+slope' baseVal
+ t_a_742 baseVal 't_a_742+slope' peakVal
+ t_a_743 peakVal 't_a_743+slope' baseVal
+ t_a_744 baseVal 't_a_744+slope' peakVal
+ t_a_745 peakVal 't_a_745+slope' baseVal
+ t_a_746 baseVal 't_a_746+slope' peakVal
+ t_a_747 peakVal 't_a_747+slope' baseVal
+ t_a_748 baseVal 't_a_748+slope' peakVal
+ t_a_749 peakVal 't_a_749+slope' baseVal
+ t_a_750 baseVal 't_a_750+slope' peakVal
+ t_a_751 peakVal 't_a_751+slope' baseVal
+ t_a_752 baseVal 't_a_752+slope' peakVal
+ t_a_753 peakVal 't_a_753+slope' baseVal
+ t_a_754 baseVal 't_a_754+slope' peakVal
+ t_a_755 peakVal 't_a_755+slope' baseVal
+ t_a_756 baseVal 't_a_756+slope' peakVal
+ t_a_757 peakVal 't_a_757+slope' baseVal
+ t_a_758 baseVal 't_a_758+slope' peakVal
+ t_a_759 peakVal 't_a_759+slope' baseVal
+ t_a_760 baseVal 't_a_760+slope' peakVal
+ t_a_761 peakVal 't_a_761+slope' baseVal
+ t_a_762 baseVal 't_a_762+slope' peakVal
+ t_a_763 peakVal 't_a_763+slope' baseVal
+ t_a_764 baseVal 't_a_764+slope' peakVal
+ t_a_765 peakVal 't_a_765+slope' baseVal
+ t_a_766 baseVal 't_a_766+slope' peakVal
+ t_a_767 peakVal 't_a_767+slope' baseVal
+ t_a_768 baseVal 't_a_768+slope' peakVal
+ t_a_769 peakVal 't_a_769+slope' baseVal
+ t_a_770 baseVal 't_a_770+slope' peakVal
+ t_a_771 peakVal 't_a_771+slope' baseVal
+ t_a_772 baseVal 't_a_772+slope' peakVal
+ t_a_773 peakVal 't_a_773+slope' baseVal
+ t_a_774 baseVal 't_a_774+slope' peakVal
+ t_a_775 peakVal 't_a_775+slope' baseVal
+ t_a_776 baseVal 't_a_776+slope' peakVal
+ t_a_777 peakVal 't_a_777+slope' baseVal
+ t_a_778 baseVal 't_a_778+slope' peakVal
+ t_a_779 peakVal 't_a_779+slope' baseVal
+ t_a_780 baseVal 't_a_780+slope' peakVal
+ t_a_781 peakVal 't_a_781+slope' baseVal
+ t_a_782 baseVal 't_a_782+slope' peakVal
+ t_a_783 peakVal 't_a_783+slope' baseVal
+ t_a_784 baseVal 't_a_784+slope' peakVal
+ t_a_785 peakVal 't_a_785+slope' baseVal
+ t_a_786 baseVal 't_a_786+slope' peakVal
+ t_a_787 peakVal 't_a_787+slope' baseVal
+ t_a_788 baseVal 't_a_788+slope' peakVal
+ t_a_789 peakVal 't_a_789+slope' baseVal
+ t_a_790 baseVal 't_a_790+slope' peakVal
+ t_a_791 peakVal 't_a_791+slope' baseVal
+ t_a_792 baseVal 't_a_792+slope' peakVal
+ t_a_793 peakVal 't_a_793+slope' baseVal
+ t_a_794 baseVal 't_a_794+slope' peakVal
+ t_a_795 peakVal 't_a_795+slope' baseVal
+ t_a_796 baseVal 't_a_796+slope' peakVal
+ t_a_797 peakVal 't_a_797+slope' baseVal
+ t_a_798 baseVal 't_a_798+slope' peakVal
+ t_a_799 peakVal 't_a_799+slope' baseVal



VINB Input_B GND PWL 0ns baseVal t_init0 baseVal 't_init0+slope' peakVal t_init1 peakVal 't_init1+slope' baseVal
+ t_b_0 baseVal 't_b_0+slope' peakVal
+ t_b_1 peakVal 't_b_1+slope' baseVal
+ t_b_2 baseVal 't_b_2+slope' peakVal
+ t_b_3 peakVal 't_b_3+slope' baseVal
+ t_b_4 baseVal 't_b_4+slope' peakVal
+ t_b_5 peakVal 't_b_5+slope' baseVal
+ t_b_6 baseVal 't_b_6+slope' peakVal
+ t_b_7 peakVal 't_b_7+slope' baseVal
+ t_b_8 baseVal 't_b_8+slope' peakVal
+ t_b_9 peakVal 't_b_9+slope' baseVal
+ t_b_10 baseVal 't_b_10+slope' peakVal
+ t_b_11 peakVal 't_b_11+slope' baseVal
+ t_b_12 baseVal 't_b_12+slope' peakVal
+ t_b_13 peakVal 't_b_13+slope' baseVal
+ t_b_14 baseVal 't_b_14+slope' peakVal
+ t_b_15 peakVal 't_b_15+slope' baseVal
+ t_b_16 baseVal 't_b_16+slope' peakVal
+ t_b_17 peakVal 't_b_17+slope' baseVal
+ t_b_18 baseVal 't_b_18+slope' peakVal
+ t_b_19 peakVal 't_b_19+slope' baseVal
+ t_b_20 baseVal 't_b_20+slope' peakVal
+ t_b_21 peakVal 't_b_21+slope' baseVal
+ t_b_22 baseVal 't_b_22+slope' peakVal
+ t_b_23 peakVal 't_b_23+slope' baseVal
+ t_b_24 baseVal 't_b_24+slope' peakVal
+ t_b_25 peakVal 't_b_25+slope' baseVal
+ t_b_26 baseVal 't_b_26+slope' peakVal
+ t_b_27 peakVal 't_b_27+slope' baseVal
+ t_b_28 baseVal 't_b_28+slope' peakVal
+ t_b_29 peakVal 't_b_29+slope' baseVal
+ t_b_30 baseVal 't_b_30+slope' peakVal
+ t_b_31 peakVal 't_b_31+slope' baseVal
+ t_b_32 baseVal 't_b_32+slope' peakVal
+ t_b_33 peakVal 't_b_33+slope' baseVal
+ t_b_34 baseVal 't_b_34+slope' peakVal
+ t_b_35 peakVal 't_b_35+slope' baseVal
+ t_b_36 baseVal 't_b_36+slope' peakVal
+ t_b_37 peakVal 't_b_37+slope' baseVal
+ t_b_38 baseVal 't_b_38+slope' peakVal
+ t_b_39 peakVal 't_b_39+slope' baseVal
+ t_b_40 baseVal 't_b_40+slope' peakVal
+ t_b_41 peakVal 't_b_41+slope' baseVal
+ t_b_42 baseVal 't_b_42+slope' peakVal
+ t_b_43 peakVal 't_b_43+slope' baseVal
+ t_b_44 baseVal 't_b_44+slope' peakVal
+ t_b_45 peakVal 't_b_45+slope' baseVal
+ t_b_46 baseVal 't_b_46+slope' peakVal
+ t_b_47 peakVal 't_b_47+slope' baseVal
+ t_b_48 baseVal 't_b_48+slope' peakVal
+ t_b_49 peakVal 't_b_49+slope' baseVal
+ t_b_50 baseVal 't_b_50+slope' peakVal
+ t_b_51 peakVal 't_b_51+slope' baseVal
+ t_b_52 baseVal 't_b_52+slope' peakVal
+ t_b_53 peakVal 't_b_53+slope' baseVal
+ t_b_54 baseVal 't_b_54+slope' peakVal
+ t_b_55 peakVal 't_b_55+slope' baseVal
+ t_b_56 baseVal 't_b_56+slope' peakVal
+ t_b_57 peakVal 't_b_57+slope' baseVal
+ t_b_58 baseVal 't_b_58+slope' peakVal
+ t_b_59 peakVal 't_b_59+slope' baseVal
+ t_b_60 baseVal 't_b_60+slope' peakVal
+ t_b_61 peakVal 't_b_61+slope' baseVal
+ t_b_62 baseVal 't_b_62+slope' peakVal
+ t_b_63 peakVal 't_b_63+slope' baseVal
+ t_b_64 baseVal 't_b_64+slope' peakVal
+ t_b_65 peakVal 't_b_65+slope' baseVal
+ t_b_66 baseVal 't_b_66+slope' peakVal
+ t_b_67 peakVal 't_b_67+slope' baseVal
+ t_b_68 baseVal 't_b_68+slope' peakVal
+ t_b_69 peakVal 't_b_69+slope' baseVal
+ t_b_70 baseVal 't_b_70+slope' peakVal
+ t_b_71 peakVal 't_b_71+slope' baseVal
+ t_b_72 baseVal 't_b_72+slope' peakVal
+ t_b_73 peakVal 't_b_73+slope' baseVal
+ t_b_74 baseVal 't_b_74+slope' peakVal
+ t_b_75 peakVal 't_b_75+slope' baseVal
+ t_b_76 baseVal 't_b_76+slope' peakVal
+ t_b_77 peakVal 't_b_77+slope' baseVal
+ t_b_78 baseVal 't_b_78+slope' peakVal
+ t_b_79 peakVal 't_b_79+slope' baseVal
+ t_b_80 baseVal 't_b_80+slope' peakVal
+ t_b_81 peakVal 't_b_81+slope' baseVal
+ t_b_82 baseVal 't_b_82+slope' peakVal
+ t_b_83 peakVal 't_b_83+slope' baseVal
+ t_b_84 baseVal 't_b_84+slope' peakVal
+ t_b_85 peakVal 't_b_85+slope' baseVal
+ t_b_86 baseVal 't_b_86+slope' peakVal
+ t_b_87 peakVal 't_b_87+slope' baseVal
+ t_b_88 baseVal 't_b_88+slope' peakVal
+ t_b_89 peakVal 't_b_89+slope' baseVal
+ t_b_90 baseVal 't_b_90+slope' peakVal
+ t_b_91 peakVal 't_b_91+slope' baseVal
+ t_b_92 baseVal 't_b_92+slope' peakVal
+ t_b_93 peakVal 't_b_93+slope' baseVal
+ t_b_94 baseVal 't_b_94+slope' peakVal
+ t_b_95 peakVal 't_b_95+slope' baseVal
+ t_b_96 baseVal 't_b_96+slope' peakVal
+ t_b_97 peakVal 't_b_97+slope' baseVal
+ t_b_98 baseVal 't_b_98+slope' peakVal
+ t_b_99 peakVal 't_b_99+slope' baseVal
+ t_b_100 baseVal 't_b_100+slope' peakVal
+ t_b_101 peakVal 't_b_101+slope' baseVal
+ t_b_102 baseVal 't_b_102+slope' peakVal
+ t_b_103 peakVal 't_b_103+slope' baseVal
+ t_b_104 baseVal 't_b_104+slope' peakVal
+ t_b_105 peakVal 't_b_105+slope' baseVal
+ t_b_106 baseVal 't_b_106+slope' peakVal
+ t_b_107 peakVal 't_b_107+slope' baseVal
+ t_b_108 baseVal 't_b_108+slope' peakVal
+ t_b_109 peakVal 't_b_109+slope' baseVal
+ t_b_110 baseVal 't_b_110+slope' peakVal
+ t_b_111 peakVal 't_b_111+slope' baseVal
+ t_b_112 baseVal 't_b_112+slope' peakVal
+ t_b_113 peakVal 't_b_113+slope' baseVal
+ t_b_114 baseVal 't_b_114+slope' peakVal
+ t_b_115 peakVal 't_b_115+slope' baseVal
+ t_b_116 baseVal 't_b_116+slope' peakVal
+ t_b_117 peakVal 't_b_117+slope' baseVal
+ t_b_118 baseVal 't_b_118+slope' peakVal
+ t_b_119 peakVal 't_b_119+slope' baseVal
+ t_b_120 baseVal 't_b_120+slope' peakVal
+ t_b_121 peakVal 't_b_121+slope' baseVal
+ t_b_122 baseVal 't_b_122+slope' peakVal
+ t_b_123 peakVal 't_b_123+slope' baseVal
+ t_b_124 baseVal 't_b_124+slope' peakVal
+ t_b_125 peakVal 't_b_125+slope' baseVal
+ t_b_126 baseVal 't_b_126+slope' peakVal
+ t_b_127 peakVal 't_b_127+slope' baseVal
+ t_b_128 baseVal 't_b_128+slope' peakVal
+ t_b_129 peakVal 't_b_129+slope' baseVal
+ t_b_130 baseVal 't_b_130+slope' peakVal
+ t_b_131 peakVal 't_b_131+slope' baseVal
+ t_b_132 baseVal 't_b_132+slope' peakVal
+ t_b_133 peakVal 't_b_133+slope' baseVal
+ t_b_134 baseVal 't_b_134+slope' peakVal
+ t_b_135 peakVal 't_b_135+slope' baseVal
+ t_b_136 baseVal 't_b_136+slope' peakVal
+ t_b_137 peakVal 't_b_137+slope' baseVal
+ t_b_138 baseVal 't_b_138+slope' peakVal
+ t_b_139 peakVal 't_b_139+slope' baseVal
+ t_b_140 baseVal 't_b_140+slope' peakVal
+ t_b_141 peakVal 't_b_141+slope' baseVal
+ t_b_142 baseVal 't_b_142+slope' peakVal
+ t_b_143 peakVal 't_b_143+slope' baseVal
+ t_b_144 baseVal 't_b_144+slope' peakVal
+ t_b_145 peakVal 't_b_145+slope' baseVal
+ t_b_146 baseVal 't_b_146+slope' peakVal
+ t_b_147 peakVal 't_b_147+slope' baseVal
+ t_b_148 baseVal 't_b_148+slope' peakVal
+ t_b_149 peakVal 't_b_149+slope' baseVal
+ t_b_150 baseVal 't_b_150+slope' peakVal
+ t_b_151 peakVal 't_b_151+slope' baseVal
+ t_b_152 baseVal 't_b_152+slope' peakVal
+ t_b_153 peakVal 't_b_153+slope' baseVal
+ t_b_154 baseVal 't_b_154+slope' peakVal
+ t_b_155 peakVal 't_b_155+slope' baseVal
+ t_b_156 baseVal 't_b_156+slope' peakVal
+ t_b_157 peakVal 't_b_157+slope' baseVal
+ t_b_158 baseVal 't_b_158+slope' peakVal
+ t_b_159 peakVal 't_b_159+slope' baseVal
+ t_b_160 baseVal 't_b_160+slope' peakVal
+ t_b_161 peakVal 't_b_161+slope' baseVal
+ t_b_162 baseVal 't_b_162+slope' peakVal
+ t_b_163 peakVal 't_b_163+slope' baseVal
+ t_b_164 baseVal 't_b_164+slope' peakVal
+ t_b_165 peakVal 't_b_165+slope' baseVal
+ t_b_166 baseVal 't_b_166+slope' peakVal
+ t_b_167 peakVal 't_b_167+slope' baseVal
+ t_b_168 baseVal 't_b_168+slope' peakVal
+ t_b_169 peakVal 't_b_169+slope' baseVal
+ t_b_170 baseVal 't_b_170+slope' peakVal
+ t_b_171 peakVal 't_b_171+slope' baseVal
+ t_b_172 baseVal 't_b_172+slope' peakVal
+ t_b_173 peakVal 't_b_173+slope' baseVal
+ t_b_174 baseVal 't_b_174+slope' peakVal
+ t_b_175 peakVal 't_b_175+slope' baseVal
+ t_b_176 baseVal 't_b_176+slope' peakVal
+ t_b_177 peakVal 't_b_177+slope' baseVal
+ t_b_178 baseVal 't_b_178+slope' peakVal
+ t_b_179 peakVal 't_b_179+slope' baseVal
+ t_b_180 baseVal 't_b_180+slope' peakVal
+ t_b_181 peakVal 't_b_181+slope' baseVal
+ t_b_182 baseVal 't_b_182+slope' peakVal
+ t_b_183 peakVal 't_b_183+slope' baseVal
+ t_b_184 baseVal 't_b_184+slope' peakVal
+ t_b_185 peakVal 't_b_185+slope' baseVal
+ t_b_186 baseVal 't_b_186+slope' peakVal
+ t_b_187 peakVal 't_b_187+slope' baseVal
+ t_b_188 baseVal 't_b_188+slope' peakVal
+ t_b_189 peakVal 't_b_189+slope' baseVal
+ t_b_190 baseVal 't_b_190+slope' peakVal
+ t_b_191 peakVal 't_b_191+slope' baseVal
+ t_b_192 baseVal 't_b_192+slope' peakVal
+ t_b_193 peakVal 't_b_193+slope' baseVal
+ t_b_194 baseVal 't_b_194+slope' peakVal
+ t_b_195 peakVal 't_b_195+slope' baseVal
+ t_b_196 baseVal 't_b_196+slope' peakVal
+ t_b_197 peakVal 't_b_197+slope' baseVal
+ t_b_198 baseVal 't_b_198+slope' peakVal
+ t_b_199 peakVal 't_b_199+slope' baseVal
+ t_b_200 baseVal 't_b_200+slope' peakVal
+ t_b_201 peakVal 't_b_201+slope' baseVal
+ t_b_202 baseVal 't_b_202+slope' peakVal
+ t_b_203 peakVal 't_b_203+slope' baseVal
+ t_b_204 baseVal 't_b_204+slope' peakVal
+ t_b_205 peakVal 't_b_205+slope' baseVal
+ t_b_206 baseVal 't_b_206+slope' peakVal
+ t_b_207 peakVal 't_b_207+slope' baseVal
+ t_b_208 baseVal 't_b_208+slope' peakVal
+ t_b_209 peakVal 't_b_209+slope' baseVal
+ t_b_210 baseVal 't_b_210+slope' peakVal
+ t_b_211 peakVal 't_b_211+slope' baseVal
+ t_b_212 baseVal 't_b_212+slope' peakVal
+ t_b_213 peakVal 't_b_213+slope' baseVal
+ t_b_214 baseVal 't_b_214+slope' peakVal
+ t_b_215 peakVal 't_b_215+slope' baseVal
+ t_b_216 baseVal 't_b_216+slope' peakVal
+ t_b_217 peakVal 't_b_217+slope' baseVal
+ t_b_218 baseVal 't_b_218+slope' peakVal
+ t_b_219 peakVal 't_b_219+slope' baseVal
+ t_b_220 baseVal 't_b_220+slope' peakVal
+ t_b_221 peakVal 't_b_221+slope' baseVal
+ t_b_222 baseVal 't_b_222+slope' peakVal
+ t_b_223 peakVal 't_b_223+slope' baseVal
+ t_b_224 baseVal 't_b_224+slope' peakVal
+ t_b_225 peakVal 't_b_225+slope' baseVal
+ t_b_226 baseVal 't_b_226+slope' peakVal
+ t_b_227 peakVal 't_b_227+slope' baseVal
+ t_b_228 baseVal 't_b_228+slope' peakVal
+ t_b_229 peakVal 't_b_229+slope' baseVal
+ t_b_230 baseVal 't_b_230+slope' peakVal
+ t_b_231 peakVal 't_b_231+slope' baseVal
+ t_b_232 baseVal 't_b_232+slope' peakVal
+ t_b_233 peakVal 't_b_233+slope' baseVal
+ t_b_234 baseVal 't_b_234+slope' peakVal
+ t_b_235 peakVal 't_b_235+slope' baseVal
+ t_b_236 baseVal 't_b_236+slope' peakVal
+ t_b_237 peakVal 't_b_237+slope' baseVal
+ t_b_238 baseVal 't_b_238+slope' peakVal
+ t_b_239 peakVal 't_b_239+slope' baseVal
+ t_b_240 baseVal 't_b_240+slope' peakVal
+ t_b_241 peakVal 't_b_241+slope' baseVal
+ t_b_242 baseVal 't_b_242+slope' peakVal
+ t_b_243 peakVal 't_b_243+slope' baseVal
+ t_b_244 baseVal 't_b_244+slope' peakVal
+ t_b_245 peakVal 't_b_245+slope' baseVal
+ t_b_246 baseVal 't_b_246+slope' peakVal
+ t_b_247 peakVal 't_b_247+slope' baseVal
+ t_b_248 baseVal 't_b_248+slope' peakVal
+ t_b_249 peakVal 't_b_249+slope' baseVal
+ t_b_250 baseVal 't_b_250+slope' peakVal
+ t_b_251 peakVal 't_b_251+slope' baseVal
+ t_b_252 baseVal 't_b_252+slope' peakVal
+ t_b_253 peakVal 't_b_253+slope' baseVal
+ t_b_254 baseVal 't_b_254+slope' peakVal
+ t_b_255 peakVal 't_b_255+slope' baseVal
+ t_b_256 baseVal 't_b_256+slope' peakVal
+ t_b_257 peakVal 't_b_257+slope' baseVal
+ t_b_258 baseVal 't_b_258+slope' peakVal
+ t_b_259 peakVal 't_b_259+slope' baseVal
+ t_b_260 baseVal 't_b_260+slope' peakVal
+ t_b_261 peakVal 't_b_261+slope' baseVal
+ t_b_262 baseVal 't_b_262+slope' peakVal
+ t_b_263 peakVal 't_b_263+slope' baseVal
+ t_b_264 baseVal 't_b_264+slope' peakVal
+ t_b_265 peakVal 't_b_265+slope' baseVal
+ t_b_266 baseVal 't_b_266+slope' peakVal
+ t_b_267 peakVal 't_b_267+slope' baseVal
+ t_b_268 baseVal 't_b_268+slope' peakVal
+ t_b_269 peakVal 't_b_269+slope' baseVal
+ t_b_270 baseVal 't_b_270+slope' peakVal
+ t_b_271 peakVal 't_b_271+slope' baseVal
+ t_b_272 baseVal 't_b_272+slope' peakVal
+ t_b_273 peakVal 't_b_273+slope' baseVal
+ t_b_274 baseVal 't_b_274+slope' peakVal
+ t_b_275 peakVal 't_b_275+slope' baseVal
+ t_b_276 baseVal 't_b_276+slope' peakVal
+ t_b_277 peakVal 't_b_277+slope' baseVal
+ t_b_278 baseVal 't_b_278+slope' peakVal
+ t_b_279 peakVal 't_b_279+slope' baseVal
+ t_b_280 baseVal 't_b_280+slope' peakVal
+ t_b_281 peakVal 't_b_281+slope' baseVal
+ t_b_282 baseVal 't_b_282+slope' peakVal
+ t_b_283 peakVal 't_b_283+slope' baseVal
+ t_b_284 baseVal 't_b_284+slope' peakVal
+ t_b_285 peakVal 't_b_285+slope' baseVal
+ t_b_286 baseVal 't_b_286+slope' peakVal
+ t_b_287 peakVal 't_b_287+slope' baseVal
+ t_b_288 baseVal 't_b_288+slope' peakVal
+ t_b_289 peakVal 't_b_289+slope' baseVal
+ t_b_290 baseVal 't_b_290+slope' peakVal
+ t_b_291 peakVal 't_b_291+slope' baseVal
+ t_b_292 baseVal 't_b_292+slope' peakVal
+ t_b_293 peakVal 't_b_293+slope' baseVal
+ t_b_294 baseVal 't_b_294+slope' peakVal
+ t_b_295 peakVal 't_b_295+slope' baseVal
+ t_b_296 baseVal 't_b_296+slope' peakVal
+ t_b_297 peakVal 't_b_297+slope' baseVal
+ t_b_298 baseVal 't_b_298+slope' peakVal
+ t_b_299 peakVal 't_b_299+slope' baseVal
+ t_b_300 baseVal 't_b_300+slope' peakVal
+ t_b_301 peakVal 't_b_301+slope' baseVal
+ t_b_302 baseVal 't_b_302+slope' peakVal
+ t_b_303 peakVal 't_b_303+slope' baseVal
+ t_b_304 baseVal 't_b_304+slope' peakVal
+ t_b_305 peakVal 't_b_305+slope' baseVal
+ t_b_306 baseVal 't_b_306+slope' peakVal
+ t_b_307 peakVal 't_b_307+slope' baseVal
+ t_b_308 baseVal 't_b_308+slope' peakVal
+ t_b_309 peakVal 't_b_309+slope' baseVal
+ t_b_310 baseVal 't_b_310+slope' peakVal
+ t_b_311 peakVal 't_b_311+slope' baseVal
+ t_b_312 baseVal 't_b_312+slope' peakVal
+ t_b_313 peakVal 't_b_313+slope' baseVal
+ t_b_314 baseVal 't_b_314+slope' peakVal
+ t_b_315 peakVal 't_b_315+slope' baseVal
+ t_b_316 baseVal 't_b_316+slope' peakVal
+ t_b_317 peakVal 't_b_317+slope' baseVal
+ t_b_318 baseVal 't_b_318+slope' peakVal
+ t_b_319 peakVal 't_b_319+slope' baseVal
+ t_b_320 baseVal 't_b_320+slope' peakVal
+ t_b_321 peakVal 't_b_321+slope' baseVal
+ t_b_322 baseVal 't_b_322+slope' peakVal
+ t_b_323 peakVal 't_b_323+slope' baseVal
+ t_b_324 baseVal 't_b_324+slope' peakVal
+ t_b_325 peakVal 't_b_325+slope' baseVal
+ t_b_326 baseVal 't_b_326+slope' peakVal
+ t_b_327 peakVal 't_b_327+slope' baseVal
+ t_b_328 baseVal 't_b_328+slope' peakVal
+ t_b_329 peakVal 't_b_329+slope' baseVal
+ t_b_330 baseVal 't_b_330+slope' peakVal
+ t_b_331 peakVal 't_b_331+slope' baseVal
+ t_b_332 baseVal 't_b_332+slope' peakVal
+ t_b_333 peakVal 't_b_333+slope' baseVal
+ t_b_334 baseVal 't_b_334+slope' peakVal
+ t_b_335 peakVal 't_b_335+slope' baseVal
+ t_b_336 baseVal 't_b_336+slope' peakVal
+ t_b_337 peakVal 't_b_337+slope' baseVal
+ t_b_338 baseVal 't_b_338+slope' peakVal
+ t_b_339 peakVal 't_b_339+slope' baseVal
+ t_b_340 baseVal 't_b_340+slope' peakVal
+ t_b_341 peakVal 't_b_341+slope' baseVal
+ t_b_342 baseVal 't_b_342+slope' peakVal
+ t_b_343 peakVal 't_b_343+slope' baseVal
+ t_b_344 baseVal 't_b_344+slope' peakVal
+ t_b_345 peakVal 't_b_345+slope' baseVal
+ t_b_346 baseVal 't_b_346+slope' peakVal
+ t_b_347 peakVal 't_b_347+slope' baseVal
+ t_b_348 baseVal 't_b_348+slope' peakVal
+ t_b_349 peakVal 't_b_349+slope' baseVal
+ t_b_350 baseVal 't_b_350+slope' peakVal
+ t_b_351 peakVal 't_b_351+slope' baseVal
+ t_b_352 baseVal 't_b_352+slope' peakVal
+ t_b_353 peakVal 't_b_353+slope' baseVal
+ t_b_354 baseVal 't_b_354+slope' peakVal
+ t_b_355 peakVal 't_b_355+slope' baseVal
+ t_b_356 baseVal 't_b_356+slope' peakVal
+ t_b_357 peakVal 't_b_357+slope' baseVal
+ t_b_358 baseVal 't_b_358+slope' peakVal
+ t_b_359 peakVal 't_b_359+slope' baseVal
+ t_b_360 baseVal 't_b_360+slope' peakVal
+ t_b_361 peakVal 't_b_361+slope' baseVal
+ t_b_362 baseVal 't_b_362+slope' peakVal
+ t_b_363 peakVal 't_b_363+slope' baseVal
+ t_b_364 baseVal 't_b_364+slope' peakVal
+ t_b_365 peakVal 't_b_365+slope' baseVal
+ t_b_366 baseVal 't_b_366+slope' peakVal
+ t_b_367 peakVal 't_b_367+slope' baseVal
+ t_b_368 baseVal 't_b_368+slope' peakVal
+ t_b_369 peakVal 't_b_369+slope' baseVal
+ t_b_370 baseVal 't_b_370+slope' peakVal
+ t_b_371 peakVal 't_b_371+slope' baseVal
+ t_b_372 baseVal 't_b_372+slope' peakVal
+ t_b_373 peakVal 't_b_373+slope' baseVal
+ t_b_374 baseVal 't_b_374+slope' peakVal
+ t_b_375 peakVal 't_b_375+slope' baseVal
+ t_b_376 baseVal 't_b_376+slope' peakVal
+ t_b_377 peakVal 't_b_377+slope' baseVal
+ t_b_378 baseVal 't_b_378+slope' peakVal
+ t_b_379 peakVal 't_b_379+slope' baseVal
+ t_b_380 baseVal 't_b_380+slope' peakVal
+ t_b_381 peakVal 't_b_381+slope' baseVal
+ t_b_382 baseVal 't_b_382+slope' peakVal
+ t_b_383 peakVal 't_b_383+slope' baseVal
+ t_b_384 baseVal 't_b_384+slope' peakVal
+ t_b_385 peakVal 't_b_385+slope' baseVal
+ t_b_386 baseVal 't_b_386+slope' peakVal
+ t_b_387 peakVal 't_b_387+slope' baseVal
+ t_b_388 baseVal 't_b_388+slope' peakVal
+ t_b_389 peakVal 't_b_389+slope' baseVal
+ t_b_390 baseVal 't_b_390+slope' peakVal
+ t_b_391 peakVal 't_b_391+slope' baseVal
+ t_b_392 baseVal 't_b_392+slope' peakVal
+ t_b_393 peakVal 't_b_393+slope' baseVal
+ t_b_394 baseVal 't_b_394+slope' peakVal
+ t_b_395 peakVal 't_b_395+slope' baseVal
+ t_b_396 baseVal 't_b_396+slope' peakVal
+ t_b_397 peakVal 't_b_397+slope' baseVal
+ t_b_398 baseVal 't_b_398+slope' peakVal
+ t_b_399 peakVal 't_b_399+slope' baseVal
+ t_b_400 baseVal 't_b_400+slope' peakVal
+ t_b_401 peakVal 't_b_401+slope' baseVal
+ t_b_402 baseVal 't_b_402+slope' peakVal
+ t_b_403 peakVal 't_b_403+slope' baseVal
+ t_b_404 baseVal 't_b_404+slope' peakVal
+ t_b_405 peakVal 't_b_405+slope' baseVal
+ t_b_406 baseVal 't_b_406+slope' peakVal
+ t_b_407 peakVal 't_b_407+slope' baseVal
+ t_b_408 baseVal 't_b_408+slope' peakVal
+ t_b_409 peakVal 't_b_409+slope' baseVal
+ t_b_410 baseVal 't_b_410+slope' peakVal
+ t_b_411 peakVal 't_b_411+slope' baseVal
+ t_b_412 baseVal 't_b_412+slope' peakVal
+ t_b_413 peakVal 't_b_413+slope' baseVal
+ t_b_414 baseVal 't_b_414+slope' peakVal
+ t_b_415 peakVal 't_b_415+slope' baseVal
+ t_b_416 baseVal 't_b_416+slope' peakVal
+ t_b_417 peakVal 't_b_417+slope' baseVal
+ t_b_418 baseVal 't_b_418+slope' peakVal
+ t_b_419 peakVal 't_b_419+slope' baseVal
+ t_b_420 baseVal 't_b_420+slope' peakVal
+ t_b_421 peakVal 't_b_421+slope' baseVal
+ t_b_422 baseVal 't_b_422+slope' peakVal
+ t_b_423 peakVal 't_b_423+slope' baseVal
+ t_b_424 baseVal 't_b_424+slope' peakVal
+ t_b_425 peakVal 't_b_425+slope' baseVal
+ t_b_426 baseVal 't_b_426+slope' peakVal
+ t_b_427 peakVal 't_b_427+slope' baseVal
+ t_b_428 baseVal 't_b_428+slope' peakVal
+ t_b_429 peakVal 't_b_429+slope' baseVal
+ t_b_430 baseVal 't_b_430+slope' peakVal
+ t_b_431 peakVal 't_b_431+slope' baseVal
+ t_b_432 baseVal 't_b_432+slope' peakVal
+ t_b_433 peakVal 't_b_433+slope' baseVal
+ t_b_434 baseVal 't_b_434+slope' peakVal
+ t_b_435 peakVal 't_b_435+slope' baseVal
+ t_b_436 baseVal 't_b_436+slope' peakVal
+ t_b_437 peakVal 't_b_437+slope' baseVal
+ t_b_438 baseVal 't_b_438+slope' peakVal
+ t_b_439 peakVal 't_b_439+slope' baseVal
+ t_b_440 baseVal 't_b_440+slope' peakVal
+ t_b_441 peakVal 't_b_441+slope' baseVal
+ t_b_442 baseVal 't_b_442+slope' peakVal
+ t_b_443 peakVal 't_b_443+slope' baseVal
+ t_b_444 baseVal 't_b_444+slope' peakVal
+ t_b_445 peakVal 't_b_445+slope' baseVal
+ t_b_446 baseVal 't_b_446+slope' peakVal
+ t_b_447 peakVal 't_b_447+slope' baseVal
+ t_b_448 baseVal 't_b_448+slope' peakVal
+ t_b_449 peakVal 't_b_449+slope' baseVal
+ t_b_450 baseVal 't_b_450+slope' peakVal
+ t_b_451 peakVal 't_b_451+slope' baseVal
+ t_b_452 baseVal 't_b_452+slope' peakVal
+ t_b_453 peakVal 't_b_453+slope' baseVal
+ t_b_454 baseVal 't_b_454+slope' peakVal
+ t_b_455 peakVal 't_b_455+slope' baseVal
+ t_b_456 baseVal 't_b_456+slope' peakVal
+ t_b_457 peakVal 't_b_457+slope' baseVal
+ t_b_458 baseVal 't_b_458+slope' peakVal
+ t_b_459 peakVal 't_b_459+slope' baseVal
+ t_b_460 baseVal 't_b_460+slope' peakVal
+ t_b_461 peakVal 't_b_461+slope' baseVal
+ t_b_462 baseVal 't_b_462+slope' peakVal
+ t_b_463 peakVal 't_b_463+slope' baseVal
+ t_b_464 baseVal 't_b_464+slope' peakVal
+ t_b_465 peakVal 't_b_465+slope' baseVal
+ t_b_466 baseVal 't_b_466+slope' peakVal
+ t_b_467 peakVal 't_b_467+slope' baseVal
+ t_b_468 baseVal 't_b_468+slope' peakVal
+ t_b_469 peakVal 't_b_469+slope' baseVal
+ t_b_470 baseVal 't_b_470+slope' peakVal
+ t_b_471 peakVal 't_b_471+slope' baseVal
+ t_b_472 baseVal 't_b_472+slope' peakVal
+ t_b_473 peakVal 't_b_473+slope' baseVal
+ t_b_474 baseVal 't_b_474+slope' peakVal
+ t_b_475 peakVal 't_b_475+slope' baseVal
+ t_b_476 baseVal 't_b_476+slope' peakVal
+ t_b_477 peakVal 't_b_477+slope' baseVal
+ t_b_478 baseVal 't_b_478+slope' peakVal
+ t_b_479 peakVal 't_b_479+slope' baseVal
+ t_b_480 baseVal 't_b_480+slope' peakVal
+ t_b_481 peakVal 't_b_481+slope' baseVal
+ t_b_482 baseVal 't_b_482+slope' peakVal
+ t_b_483 peakVal 't_b_483+slope' baseVal
+ t_b_484 baseVal 't_b_484+slope' peakVal
+ t_b_485 peakVal 't_b_485+slope' baseVal
+ t_b_486 baseVal 't_b_486+slope' peakVal
+ t_b_487 peakVal 't_b_487+slope' baseVal
+ t_b_488 baseVal 't_b_488+slope' peakVal
+ t_b_489 peakVal 't_b_489+slope' baseVal
+ t_b_490 baseVal 't_b_490+slope' peakVal
+ t_b_491 peakVal 't_b_491+slope' baseVal
+ t_b_492 baseVal 't_b_492+slope' peakVal
+ t_b_493 peakVal 't_b_493+slope' baseVal
+ t_b_494 baseVal 't_b_494+slope' peakVal
+ t_b_495 peakVal 't_b_495+slope' baseVal
+ t_b_496 baseVal 't_b_496+slope' peakVal
+ t_b_497 peakVal 't_b_497+slope' baseVal
+ t_b_498 baseVal 't_b_498+slope' peakVal
+ t_b_499 peakVal 't_b_499+slope' baseVal
+ t_b_500 baseVal 't_b_500+slope' peakVal
+ t_b_501 peakVal 't_b_501+slope' baseVal
+ t_b_502 baseVal 't_b_502+slope' peakVal
+ t_b_503 peakVal 't_b_503+slope' baseVal
+ t_b_504 baseVal 't_b_504+slope' peakVal
+ t_b_505 peakVal 't_b_505+slope' baseVal
+ t_b_506 baseVal 't_b_506+slope' peakVal
+ t_b_507 peakVal 't_b_507+slope' baseVal
+ t_b_508 baseVal 't_b_508+slope' peakVal
+ t_b_509 peakVal 't_b_509+slope' baseVal
+ t_b_510 baseVal 't_b_510+slope' peakVal
+ t_b_511 peakVal 't_b_511+slope' baseVal
+ t_b_512 baseVal 't_b_512+slope' peakVal
+ t_b_513 peakVal 't_b_513+slope' baseVal
+ t_b_514 baseVal 't_b_514+slope' peakVal
+ t_b_515 peakVal 't_b_515+slope' baseVal
+ t_b_516 baseVal 't_b_516+slope' peakVal
+ t_b_517 peakVal 't_b_517+slope' baseVal
+ t_b_518 baseVal 't_b_518+slope' peakVal
+ t_b_519 peakVal 't_b_519+slope' baseVal
+ t_b_520 baseVal 't_b_520+slope' peakVal
+ t_b_521 peakVal 't_b_521+slope' baseVal
+ t_b_522 baseVal 't_b_522+slope' peakVal
+ t_b_523 peakVal 't_b_523+slope' baseVal
+ t_b_524 baseVal 't_b_524+slope' peakVal
+ t_b_525 peakVal 't_b_525+slope' baseVal
+ t_b_526 baseVal 't_b_526+slope' peakVal
+ t_b_527 peakVal 't_b_527+slope' baseVal
+ t_b_528 baseVal 't_b_528+slope' peakVal
+ t_b_529 peakVal 't_b_529+slope' baseVal
+ t_b_530 baseVal 't_b_530+slope' peakVal
+ t_b_531 peakVal 't_b_531+slope' baseVal
+ t_b_532 baseVal 't_b_532+slope' peakVal
+ t_b_533 peakVal 't_b_533+slope' baseVal
+ t_b_534 baseVal 't_b_534+slope' peakVal
+ t_b_535 peakVal 't_b_535+slope' baseVal
+ t_b_536 baseVal 't_b_536+slope' peakVal
+ t_b_537 peakVal 't_b_537+slope' baseVal
+ t_b_538 baseVal 't_b_538+slope' peakVal
+ t_b_539 peakVal 't_b_539+slope' baseVal
+ t_b_540 baseVal 't_b_540+slope' peakVal
+ t_b_541 peakVal 't_b_541+slope' baseVal
+ t_b_542 baseVal 't_b_542+slope' peakVal
+ t_b_543 peakVal 't_b_543+slope' baseVal
+ t_b_544 baseVal 't_b_544+slope' peakVal
+ t_b_545 peakVal 't_b_545+slope' baseVal
+ t_b_546 baseVal 't_b_546+slope' peakVal
+ t_b_547 peakVal 't_b_547+slope' baseVal
+ t_b_548 baseVal 't_b_548+slope' peakVal
+ t_b_549 peakVal 't_b_549+slope' baseVal
+ t_b_550 baseVal 't_b_550+slope' peakVal
+ t_b_551 peakVal 't_b_551+slope' baseVal
+ t_b_552 baseVal 't_b_552+slope' peakVal
+ t_b_553 peakVal 't_b_553+slope' baseVal
+ t_b_554 baseVal 't_b_554+slope' peakVal
+ t_b_555 peakVal 't_b_555+slope' baseVal
+ t_b_556 baseVal 't_b_556+slope' peakVal
+ t_b_557 peakVal 't_b_557+slope' baseVal
+ t_b_558 baseVal 't_b_558+slope' peakVal
+ t_b_559 peakVal 't_b_559+slope' baseVal
+ t_b_560 baseVal 't_b_560+slope' peakVal
+ t_b_561 peakVal 't_b_561+slope' baseVal
+ t_b_562 baseVal 't_b_562+slope' peakVal
+ t_b_563 peakVal 't_b_563+slope' baseVal
+ t_b_564 baseVal 't_b_564+slope' peakVal
+ t_b_565 peakVal 't_b_565+slope' baseVal
+ t_b_566 baseVal 't_b_566+slope' peakVal
+ t_b_567 peakVal 't_b_567+slope' baseVal
+ t_b_568 baseVal 't_b_568+slope' peakVal
+ t_b_569 peakVal 't_b_569+slope' baseVal
+ t_b_570 baseVal 't_b_570+slope' peakVal
+ t_b_571 peakVal 't_b_571+slope' baseVal
+ t_b_572 baseVal 't_b_572+slope' peakVal
+ t_b_573 peakVal 't_b_573+slope' baseVal
+ t_b_574 baseVal 't_b_574+slope' peakVal
+ t_b_575 peakVal 't_b_575+slope' baseVal
+ t_b_576 baseVal 't_b_576+slope' peakVal
+ t_b_577 peakVal 't_b_577+slope' baseVal
+ t_b_578 baseVal 't_b_578+slope' peakVal
+ t_b_579 peakVal 't_b_579+slope' baseVal
+ t_b_580 baseVal 't_b_580+slope' peakVal
+ t_b_581 peakVal 't_b_581+slope' baseVal
+ t_b_582 baseVal 't_b_582+slope' peakVal
+ t_b_583 peakVal 't_b_583+slope' baseVal
+ t_b_584 baseVal 't_b_584+slope' peakVal
+ t_b_585 peakVal 't_b_585+slope' baseVal
+ t_b_586 baseVal 't_b_586+slope' peakVal
+ t_b_587 peakVal 't_b_587+slope' baseVal
+ t_b_588 baseVal 't_b_588+slope' peakVal
+ t_b_589 peakVal 't_b_589+slope' baseVal
+ t_b_590 baseVal 't_b_590+slope' peakVal
+ t_b_591 peakVal 't_b_591+slope' baseVal
+ t_b_592 baseVal 't_b_592+slope' peakVal
+ t_b_593 peakVal 't_b_593+slope' baseVal
+ t_b_594 baseVal 't_b_594+slope' peakVal
+ t_b_595 peakVal 't_b_595+slope' baseVal
+ t_b_596 baseVal 't_b_596+slope' peakVal
+ t_b_597 peakVal 't_b_597+slope' baseVal
+ t_b_598 baseVal 't_b_598+slope' peakVal
+ t_b_599 peakVal 't_b_599+slope' baseVal
+ t_b_600 baseVal 't_b_600+slope' peakVal
+ t_b_601 peakVal 't_b_601+slope' baseVal
+ t_b_602 baseVal 't_b_602+slope' peakVal
+ t_b_603 peakVal 't_b_603+slope' baseVal
+ t_b_604 baseVal 't_b_604+slope' peakVal
+ t_b_605 peakVal 't_b_605+slope' baseVal
+ t_b_606 baseVal 't_b_606+slope' peakVal
+ t_b_607 peakVal 't_b_607+slope' baseVal
+ t_b_608 baseVal 't_b_608+slope' peakVal
+ t_b_609 peakVal 't_b_609+slope' baseVal
+ t_b_610 baseVal 't_b_610+slope' peakVal
+ t_b_611 peakVal 't_b_611+slope' baseVal
+ t_b_612 baseVal 't_b_612+slope' peakVal
+ t_b_613 peakVal 't_b_613+slope' baseVal
+ t_b_614 baseVal 't_b_614+slope' peakVal
+ t_b_615 peakVal 't_b_615+slope' baseVal
+ t_b_616 baseVal 't_b_616+slope' peakVal
+ t_b_617 peakVal 't_b_617+slope' baseVal
+ t_b_618 baseVal 't_b_618+slope' peakVal
+ t_b_619 peakVal 't_b_619+slope' baseVal
+ t_b_620 baseVal 't_b_620+slope' peakVal
+ t_b_621 peakVal 't_b_621+slope' baseVal
+ t_b_622 baseVal 't_b_622+slope' peakVal
+ t_b_623 peakVal 't_b_623+slope' baseVal
+ t_b_624 baseVal 't_b_624+slope' peakVal
+ t_b_625 peakVal 't_b_625+slope' baseVal
+ t_b_626 baseVal 't_b_626+slope' peakVal
+ t_b_627 peakVal 't_b_627+slope' baseVal
+ t_b_628 baseVal 't_b_628+slope' peakVal
+ t_b_629 peakVal 't_b_629+slope' baseVal
+ t_b_630 baseVal 't_b_630+slope' peakVal
+ t_b_631 peakVal 't_b_631+slope' baseVal
+ t_b_632 baseVal 't_b_632+slope' peakVal
+ t_b_633 peakVal 't_b_633+slope' baseVal
+ t_b_634 baseVal 't_b_634+slope' peakVal
+ t_b_635 peakVal 't_b_635+slope' baseVal
+ t_b_636 baseVal 't_b_636+slope' peakVal
+ t_b_637 peakVal 't_b_637+slope' baseVal
+ t_b_638 baseVal 't_b_638+slope' peakVal
+ t_b_639 peakVal 't_b_639+slope' baseVal
+ t_b_640 baseVal 't_b_640+slope' peakVal
+ t_b_641 peakVal 't_b_641+slope' baseVal
+ t_b_642 baseVal 't_b_642+slope' peakVal
+ t_b_643 peakVal 't_b_643+slope' baseVal
+ t_b_644 baseVal 't_b_644+slope' peakVal
+ t_b_645 peakVal 't_b_645+slope' baseVal
+ t_b_646 baseVal 't_b_646+slope' peakVal
+ t_b_647 peakVal 't_b_647+slope' baseVal
+ t_b_648 baseVal 't_b_648+slope' peakVal
+ t_b_649 peakVal 't_b_649+slope' baseVal
+ t_b_650 baseVal 't_b_650+slope' peakVal
+ t_b_651 peakVal 't_b_651+slope' baseVal
+ t_b_652 baseVal 't_b_652+slope' peakVal
+ t_b_653 peakVal 't_b_653+slope' baseVal
+ t_b_654 baseVal 't_b_654+slope' peakVal
+ t_b_655 peakVal 't_b_655+slope' baseVal
+ t_b_656 baseVal 't_b_656+slope' peakVal
+ t_b_657 peakVal 't_b_657+slope' baseVal
+ t_b_658 baseVal 't_b_658+slope' peakVal
+ t_b_659 peakVal 't_b_659+slope' baseVal
+ t_b_660 baseVal 't_b_660+slope' peakVal
+ t_b_661 peakVal 't_b_661+slope' baseVal
+ t_b_662 baseVal 't_b_662+slope' peakVal
+ t_b_663 peakVal 't_b_663+slope' baseVal
+ t_b_664 baseVal 't_b_664+slope' peakVal
+ t_b_665 peakVal 't_b_665+slope' baseVal
+ t_b_666 baseVal 't_b_666+slope' peakVal
+ t_b_667 peakVal 't_b_667+slope' baseVal
+ t_b_668 baseVal 't_b_668+slope' peakVal
+ t_b_669 peakVal 't_b_669+slope' baseVal
+ t_b_670 baseVal 't_b_670+slope' peakVal
+ t_b_671 peakVal 't_b_671+slope' baseVal
+ t_b_672 baseVal 't_b_672+slope' peakVal
+ t_b_673 peakVal 't_b_673+slope' baseVal
+ t_b_674 baseVal 't_b_674+slope' peakVal
+ t_b_675 peakVal 't_b_675+slope' baseVal
+ t_b_676 baseVal 't_b_676+slope' peakVal
+ t_b_677 peakVal 't_b_677+slope' baseVal
+ t_b_678 baseVal 't_b_678+slope' peakVal
+ t_b_679 peakVal 't_b_679+slope' baseVal
+ t_b_680 baseVal 't_b_680+slope' peakVal
+ t_b_681 peakVal 't_b_681+slope' baseVal
+ t_b_682 baseVal 't_b_682+slope' peakVal
+ t_b_683 peakVal 't_b_683+slope' baseVal
+ t_b_684 baseVal 't_b_684+slope' peakVal
+ t_b_685 peakVal 't_b_685+slope' baseVal
+ t_b_686 baseVal 't_b_686+slope' peakVal
+ t_b_687 peakVal 't_b_687+slope' baseVal
+ t_b_688 baseVal 't_b_688+slope' peakVal
+ t_b_689 peakVal 't_b_689+slope' baseVal
+ t_b_690 baseVal 't_b_690+slope' peakVal
+ t_b_691 peakVal 't_b_691+slope' baseVal
+ t_b_692 baseVal 't_b_692+slope' peakVal
+ t_b_693 peakVal 't_b_693+slope' baseVal
+ t_b_694 baseVal 't_b_694+slope' peakVal
+ t_b_695 peakVal 't_b_695+slope' baseVal
+ t_b_696 baseVal 't_b_696+slope' peakVal
+ t_b_697 peakVal 't_b_697+slope' baseVal
+ t_b_698 baseVal 't_b_698+slope' peakVal
+ t_b_699 peakVal 't_b_699+slope' baseVal
+ t_b_700 baseVal 't_b_700+slope' peakVal
+ t_b_701 peakVal 't_b_701+slope' baseVal
+ t_b_702 baseVal 't_b_702+slope' peakVal
+ t_b_703 peakVal 't_b_703+slope' baseVal
+ t_b_704 baseVal 't_b_704+slope' peakVal
+ t_b_705 peakVal 't_b_705+slope' baseVal
+ t_b_706 baseVal 't_b_706+slope' peakVal
+ t_b_707 peakVal 't_b_707+slope' baseVal
+ t_b_708 baseVal 't_b_708+slope' peakVal
+ t_b_709 peakVal 't_b_709+slope' baseVal
+ t_b_710 baseVal 't_b_710+slope' peakVal
+ t_b_711 peakVal 't_b_711+slope' baseVal
+ t_b_712 baseVal 't_b_712+slope' peakVal
+ t_b_713 peakVal 't_b_713+slope' baseVal
+ t_b_714 baseVal 't_b_714+slope' peakVal
+ t_b_715 peakVal 't_b_715+slope' baseVal
+ t_b_716 baseVal 't_b_716+slope' peakVal
+ t_b_717 peakVal 't_b_717+slope' baseVal
+ t_b_718 baseVal 't_b_718+slope' peakVal
+ t_b_719 peakVal 't_b_719+slope' baseVal
+ t_b_720 baseVal 't_b_720+slope' peakVal
+ t_b_721 peakVal 't_b_721+slope' baseVal
+ t_b_722 baseVal 't_b_722+slope' peakVal
+ t_b_723 peakVal 't_b_723+slope' baseVal
+ t_b_724 baseVal 't_b_724+slope' peakVal
+ t_b_725 peakVal 't_b_725+slope' baseVal
+ t_b_726 baseVal 't_b_726+slope' peakVal
+ t_b_727 peakVal 't_b_727+slope' baseVal
+ t_b_728 baseVal 't_b_728+slope' peakVal
+ t_b_729 peakVal 't_b_729+slope' baseVal
+ t_b_730 baseVal 't_b_730+slope' peakVal
+ t_b_731 peakVal 't_b_731+slope' baseVal
+ t_b_732 baseVal 't_b_732+slope' peakVal
+ t_b_733 peakVal 't_b_733+slope' baseVal
+ t_b_734 baseVal 't_b_734+slope' peakVal
+ t_b_735 peakVal 't_b_735+slope' baseVal
+ t_b_736 baseVal 't_b_736+slope' peakVal
+ t_b_737 peakVal 't_b_737+slope' baseVal
+ t_b_738 baseVal 't_b_738+slope' peakVal
+ t_b_739 peakVal 't_b_739+slope' baseVal
+ t_b_740 baseVal 't_b_740+slope' peakVal
+ t_b_741 peakVal 't_b_741+slope' baseVal
+ t_b_742 baseVal 't_b_742+slope' peakVal
+ t_b_743 peakVal 't_b_743+slope' baseVal
+ t_b_744 baseVal 't_b_744+slope' peakVal
+ t_b_745 peakVal 't_b_745+slope' baseVal
+ t_b_746 baseVal 't_b_746+slope' peakVal
+ t_b_747 peakVal 't_b_747+slope' baseVal
+ t_b_748 baseVal 't_b_748+slope' peakVal
+ t_b_749 peakVal 't_b_749+slope' baseVal
+ t_b_750 baseVal 't_b_750+slope' peakVal
+ t_b_751 peakVal 't_b_751+slope' baseVal
+ t_b_752 baseVal 't_b_752+slope' peakVal
+ t_b_753 peakVal 't_b_753+slope' baseVal
+ t_b_754 baseVal 't_b_754+slope' peakVal
+ t_b_755 peakVal 't_b_755+slope' baseVal
+ t_b_756 baseVal 't_b_756+slope' peakVal
+ t_b_757 peakVal 't_b_757+slope' baseVal
+ t_b_758 baseVal 't_b_758+slope' peakVal
+ t_b_759 peakVal 't_b_759+slope' baseVal
+ t_b_760 baseVal 't_b_760+slope' peakVal
+ t_b_761 peakVal 't_b_761+slope' baseVal
+ t_b_762 baseVal 't_b_762+slope' peakVal
+ t_b_763 peakVal 't_b_763+slope' baseVal
+ t_b_764 baseVal 't_b_764+slope' peakVal
+ t_b_765 peakVal 't_b_765+slope' baseVal
+ t_b_766 baseVal 't_b_766+slope' peakVal
+ t_b_767 peakVal 't_b_767+slope' baseVal
+ t_b_768 baseVal 't_b_768+slope' peakVal
+ t_b_769 peakVal 't_b_769+slope' baseVal
+ t_b_770 baseVal 't_b_770+slope' peakVal
+ t_b_771 peakVal 't_b_771+slope' baseVal
+ t_b_772 baseVal 't_b_772+slope' peakVal
+ t_b_773 peakVal 't_b_773+slope' baseVal
+ t_b_774 baseVal 't_b_774+slope' peakVal
+ t_b_775 peakVal 't_b_775+slope' baseVal
+ t_b_776 baseVal 't_b_776+slope' peakVal
+ t_b_777 peakVal 't_b_777+slope' baseVal
+ t_b_778 baseVal 't_b_778+slope' peakVal
+ t_b_779 peakVal 't_b_779+slope' baseVal
+ t_b_780 baseVal 't_b_780+slope' peakVal
+ t_b_781 peakVal 't_b_781+slope' baseVal
+ t_b_782 baseVal 't_b_782+slope' peakVal
+ t_b_783 peakVal 't_b_783+slope' baseVal
+ t_b_784 baseVal 't_b_784+slope' peakVal
+ t_b_785 peakVal 't_b_785+slope' baseVal
+ t_b_786 baseVal 't_b_786+slope' peakVal
+ t_b_787 peakVal 't_b_787+slope' baseVal
+ t_b_788 baseVal 't_b_788+slope' peakVal
+ t_b_789 peakVal 't_b_789+slope' baseVal
+ t_b_790 baseVal 't_b_790+slope' peakVal
+ t_b_791 peakVal 't_b_791+slope' baseVal
+ t_b_792 baseVal 't_b_792+slope' peakVal
+ t_b_793 peakVal 't_b_793+slope' baseVal
+ t_b_794 baseVal 't_b_794+slope' peakVal
+ t_b_795 peakVal 't_b_795+slope' baseVal
+ t_b_796 baseVal 't_b_796+slope' peakVal
+ t_b_797 peakVal 't_b_797+slope' baseVal
+ t_b_798 baseVal 't_b_798+slope' peakVal
+ t_b_799 peakVal 't_b_799+slope' baseVal



*circuit

XBUFFER_A Input_A A VDD VDD GND GND BUF_X8
XBUFFER_B Input_B B VDD VDD GND GND BUF_X8
XCGATE A B Z VDD VDD GND GND CGATE
XBUFFER_Z Z Output VDD VDD GND GND BUF_X8
C_TERM Output GND 0.0779pF

.PROBE TRAN V(A) V(B) V(Z)
.TRAN 0.1ps tend
.END
module parallel_NOR_chains_50_stages(IN_A1, IN_A2, OUT_Z1, OUT_Z2);
       input IN_A1, IN_A2;
       output OUT_Z1, OUT_Z2;


       wire STAGE_0_OUT_1, STAGE_0_OUT_2;
       NOR2_X2 X_NOR_STAGE_0_1 (.A1(IN_A1), .A2(IN_A2), .ZN(STAGE_0_OUT_1));
       NOR2_X2 X_NOR_STAGE_0_2 (.A1(IN_A1), .A2(IN_A2), .ZN(STAGE_0_OUT_2));

       wire STAGE_1_OUT_1, STAGE_1_OUT_2;
       NOR2_X2 X_NOR_STAGE_1_1 (.A1(STAGE_0_OUT_1), .A2(STAGE_0_OUT_2), .ZN(STAGE_1_OUT_1));
       NOR2_X2 X_NOR_STAGE_1_2 (.A1(STAGE_0_OUT_1), .A2(STAGE_0_OUT_2), .ZN(STAGE_1_OUT_2));

       wire STAGE_2_OUT_1, STAGE_2_OUT_2;
       NOR2_X2 X_NOR_STAGE_2_1 (.A1(STAGE_1_OUT_1), .A2(STAGE_1_OUT_2), .ZN(STAGE_2_OUT_1));
       NOR2_X2 X_NOR_STAGE_2_2 (.A1(STAGE_1_OUT_1), .A2(STAGE_1_OUT_2), .ZN(STAGE_2_OUT_2));

       wire STAGE_3_OUT_1, STAGE_3_OUT_2;
       NOR2_X2 X_NOR_STAGE_3_1 (.A1(STAGE_2_OUT_1), .A2(STAGE_2_OUT_2), .ZN(STAGE_3_OUT_1));
       NOR2_X2 X_NOR_STAGE_3_2 (.A1(STAGE_2_OUT_1), .A2(STAGE_2_OUT_2), .ZN(STAGE_3_OUT_2));

       wire STAGE_4_OUT_1, STAGE_4_OUT_2;
       NOR2_X2 X_NOR_STAGE_4_1 (.A1(STAGE_3_OUT_1), .A2(STAGE_3_OUT_2), .ZN(STAGE_4_OUT_1));
       NOR2_X2 X_NOR_STAGE_4_2 (.A1(STAGE_3_OUT_1), .A2(STAGE_3_OUT_2), .ZN(STAGE_4_OUT_2));

       wire STAGE_5_OUT_1, STAGE_5_OUT_2;
       NOR2_X2 X_NOR_STAGE_5_1 (.A1(STAGE_4_OUT_1), .A2(STAGE_4_OUT_2), .ZN(STAGE_5_OUT_1));
       NOR2_X2 X_NOR_STAGE_5_2 (.A1(STAGE_4_OUT_1), .A2(STAGE_4_OUT_2), .ZN(STAGE_5_OUT_2));

       wire STAGE_6_OUT_1, STAGE_6_OUT_2;
       NOR2_X2 X_NOR_STAGE_6_1 (.A1(STAGE_5_OUT_1), .A2(STAGE_5_OUT_2), .ZN(STAGE_6_OUT_1));
       NOR2_X2 X_NOR_STAGE_6_2 (.A1(STAGE_5_OUT_1), .A2(STAGE_5_OUT_2), .ZN(STAGE_6_OUT_2));

       wire STAGE_7_OUT_1, STAGE_7_OUT_2;
       NOR2_X2 X_NOR_STAGE_7_1 (.A1(STAGE_6_OUT_1), .A2(STAGE_6_OUT_2), .ZN(STAGE_7_OUT_1));
       NOR2_X2 X_NOR_STAGE_7_2 (.A1(STAGE_6_OUT_1), .A2(STAGE_6_OUT_2), .ZN(STAGE_7_OUT_2));

       wire STAGE_8_OUT_1, STAGE_8_OUT_2;
       NOR2_X2 X_NOR_STAGE_8_1 (.A1(STAGE_7_OUT_1), .A2(STAGE_7_OUT_2), .ZN(STAGE_8_OUT_1));
       NOR2_X2 X_NOR_STAGE_8_2 (.A1(STAGE_7_OUT_1), .A2(STAGE_7_OUT_2), .ZN(STAGE_8_OUT_2));

       wire STAGE_9_OUT_1, STAGE_9_OUT_2;
       NOR2_X2 X_NOR_STAGE_9_1 (.A1(STAGE_8_OUT_1), .A2(STAGE_8_OUT_2), .ZN(STAGE_9_OUT_1));
       NOR2_X2 X_NOR_STAGE_9_2 (.A1(STAGE_8_OUT_1), .A2(STAGE_8_OUT_2), .ZN(STAGE_9_OUT_2));

       wire STAGE_10_OUT_1, STAGE_10_OUT_2;
       NOR2_X2 X_NOR_STAGE_10_1 (.A1(STAGE_9_OUT_1), .A2(STAGE_9_OUT_2), .ZN(STAGE_10_OUT_1));
       NOR2_X2 X_NOR_STAGE_10_2 (.A1(STAGE_9_OUT_1), .A2(STAGE_9_OUT_2), .ZN(STAGE_10_OUT_2));

       wire STAGE_11_OUT_1, STAGE_11_OUT_2;
       NOR2_X2 X_NOR_STAGE_11_1 (.A1(STAGE_10_OUT_1), .A2(STAGE_10_OUT_2), .ZN(STAGE_11_OUT_1));
       NOR2_X2 X_NOR_STAGE_11_2 (.A1(STAGE_10_OUT_1), .A2(STAGE_10_OUT_2), .ZN(STAGE_11_OUT_2));

       wire STAGE_12_OUT_1, STAGE_12_OUT_2;
       NOR2_X2 X_NOR_STAGE_12_1 (.A1(STAGE_11_OUT_1), .A2(STAGE_11_OUT_2), .ZN(STAGE_12_OUT_1));
       NOR2_X2 X_NOR_STAGE_12_2 (.A1(STAGE_11_OUT_1), .A2(STAGE_11_OUT_2), .ZN(STAGE_12_OUT_2));

       wire STAGE_13_OUT_1, STAGE_13_OUT_2;
       NOR2_X2 X_NOR_STAGE_13_1 (.A1(STAGE_12_OUT_1), .A2(STAGE_12_OUT_2), .ZN(STAGE_13_OUT_1));
       NOR2_X2 X_NOR_STAGE_13_2 (.A1(STAGE_12_OUT_1), .A2(STAGE_12_OUT_2), .ZN(STAGE_13_OUT_2));

       wire STAGE_14_OUT_1, STAGE_14_OUT_2;
       NOR2_X2 X_NOR_STAGE_14_1 (.A1(STAGE_13_OUT_1), .A2(STAGE_13_OUT_2), .ZN(STAGE_14_OUT_1));
       NOR2_X2 X_NOR_STAGE_14_2 (.A1(STAGE_13_OUT_1), .A2(STAGE_13_OUT_2), .ZN(STAGE_14_OUT_2));

       wire STAGE_15_OUT_1, STAGE_15_OUT_2;
       NOR2_X2 X_NOR_STAGE_15_1 (.A1(STAGE_14_OUT_1), .A2(STAGE_14_OUT_2), .ZN(STAGE_15_OUT_1));
       NOR2_X2 X_NOR_STAGE_15_2 (.A1(STAGE_14_OUT_1), .A2(STAGE_14_OUT_2), .ZN(STAGE_15_OUT_2));

       wire STAGE_16_OUT_1, STAGE_16_OUT_2;
       NOR2_X2 X_NOR_STAGE_16_1 (.A1(STAGE_15_OUT_1), .A2(STAGE_15_OUT_2), .ZN(STAGE_16_OUT_1));
       NOR2_X2 X_NOR_STAGE_16_2 (.A1(STAGE_15_OUT_1), .A2(STAGE_15_OUT_2), .ZN(STAGE_16_OUT_2));

       wire STAGE_17_OUT_1, STAGE_17_OUT_2;
       NOR2_X2 X_NOR_STAGE_17_1 (.A1(STAGE_16_OUT_1), .A2(STAGE_16_OUT_2), .ZN(STAGE_17_OUT_1));
       NOR2_X2 X_NOR_STAGE_17_2 (.A1(STAGE_16_OUT_1), .A2(STAGE_16_OUT_2), .ZN(STAGE_17_OUT_2));

       wire STAGE_18_OUT_1, STAGE_18_OUT_2;
       NOR2_X2 X_NOR_STAGE_18_1 (.A1(STAGE_17_OUT_1), .A2(STAGE_17_OUT_2), .ZN(STAGE_18_OUT_1));
       NOR2_X2 X_NOR_STAGE_18_2 (.A1(STAGE_17_OUT_1), .A2(STAGE_17_OUT_2), .ZN(STAGE_18_OUT_2));

       wire STAGE_19_OUT_1, STAGE_19_OUT_2;
       NOR2_X2 X_NOR_STAGE_19_1 (.A1(STAGE_18_OUT_1), .A2(STAGE_18_OUT_2), .ZN(STAGE_19_OUT_1));
       NOR2_X2 X_NOR_STAGE_19_2 (.A1(STAGE_18_OUT_1), .A2(STAGE_18_OUT_2), .ZN(STAGE_19_OUT_2));

       wire STAGE_20_OUT_1, STAGE_20_OUT_2;
       NOR2_X2 X_NOR_STAGE_20_1 (.A1(STAGE_19_OUT_1), .A2(STAGE_19_OUT_2), .ZN(STAGE_20_OUT_1));
       NOR2_X2 X_NOR_STAGE_20_2 (.A1(STAGE_19_OUT_1), .A2(STAGE_19_OUT_2), .ZN(STAGE_20_OUT_2));

       wire STAGE_21_OUT_1, STAGE_21_OUT_2;
       NOR2_X2 X_NOR_STAGE_21_1 (.A1(STAGE_20_OUT_1), .A2(STAGE_20_OUT_2), .ZN(STAGE_21_OUT_1));
       NOR2_X2 X_NOR_STAGE_21_2 (.A1(STAGE_20_OUT_1), .A2(STAGE_20_OUT_2), .ZN(STAGE_21_OUT_2));

       wire STAGE_22_OUT_1, STAGE_22_OUT_2;
       NOR2_X2 X_NOR_STAGE_22_1 (.A1(STAGE_21_OUT_1), .A2(STAGE_21_OUT_2), .ZN(STAGE_22_OUT_1));
       NOR2_X2 X_NOR_STAGE_22_2 (.A1(STAGE_21_OUT_1), .A2(STAGE_21_OUT_2), .ZN(STAGE_22_OUT_2));

       wire STAGE_23_OUT_1, STAGE_23_OUT_2;
       NOR2_X2 X_NOR_STAGE_23_1 (.A1(STAGE_22_OUT_1), .A2(STAGE_22_OUT_2), .ZN(STAGE_23_OUT_1));
       NOR2_X2 X_NOR_STAGE_23_2 (.A1(STAGE_22_OUT_1), .A2(STAGE_22_OUT_2), .ZN(STAGE_23_OUT_2));

       wire STAGE_24_OUT_1, STAGE_24_OUT_2;
       NOR2_X2 X_NOR_STAGE_24_1 (.A1(STAGE_23_OUT_1), .A2(STAGE_23_OUT_2), .ZN(STAGE_24_OUT_1));
       NOR2_X2 X_NOR_STAGE_24_2 (.A1(STAGE_23_OUT_1), .A2(STAGE_23_OUT_2), .ZN(STAGE_24_OUT_2));

       wire STAGE_25_OUT_1, STAGE_25_OUT_2;
       NOR2_X2 X_NOR_STAGE_25_1 (.A1(STAGE_24_OUT_1), .A2(STAGE_24_OUT_2), .ZN(STAGE_25_OUT_1));
       NOR2_X2 X_NOR_STAGE_25_2 (.A1(STAGE_24_OUT_1), .A2(STAGE_24_OUT_2), .ZN(STAGE_25_OUT_2));

       wire STAGE_26_OUT_1, STAGE_26_OUT_2;
       NOR2_X2 X_NOR_STAGE_26_1 (.A1(STAGE_25_OUT_1), .A2(STAGE_25_OUT_2), .ZN(STAGE_26_OUT_1));
       NOR2_X2 X_NOR_STAGE_26_2 (.A1(STAGE_25_OUT_1), .A2(STAGE_25_OUT_2), .ZN(STAGE_26_OUT_2));

       wire STAGE_27_OUT_1, STAGE_27_OUT_2;
       NOR2_X2 X_NOR_STAGE_27_1 (.A1(STAGE_26_OUT_1), .A2(STAGE_26_OUT_2), .ZN(STAGE_27_OUT_1));
       NOR2_X2 X_NOR_STAGE_27_2 (.A1(STAGE_26_OUT_1), .A2(STAGE_26_OUT_2), .ZN(STAGE_27_OUT_2));

       wire STAGE_28_OUT_1, STAGE_28_OUT_2;
       NOR2_X2 X_NOR_STAGE_28_1 (.A1(STAGE_27_OUT_1), .A2(STAGE_27_OUT_2), .ZN(STAGE_28_OUT_1));
       NOR2_X2 X_NOR_STAGE_28_2 (.A1(STAGE_27_OUT_1), .A2(STAGE_27_OUT_2), .ZN(STAGE_28_OUT_2));

       wire STAGE_29_OUT_1, STAGE_29_OUT_2;
       NOR2_X2 X_NOR_STAGE_29_1 (.A1(STAGE_28_OUT_1), .A2(STAGE_28_OUT_2), .ZN(STAGE_29_OUT_1));
       NOR2_X2 X_NOR_STAGE_29_2 (.A1(STAGE_28_OUT_1), .A2(STAGE_28_OUT_2), .ZN(STAGE_29_OUT_2));

       wire STAGE_30_OUT_1, STAGE_30_OUT_2;
       NOR2_X2 X_NOR_STAGE_30_1 (.A1(STAGE_29_OUT_1), .A2(STAGE_29_OUT_2), .ZN(STAGE_30_OUT_1));
       NOR2_X2 X_NOR_STAGE_30_2 (.A1(STAGE_29_OUT_1), .A2(STAGE_29_OUT_2), .ZN(STAGE_30_OUT_2));

       wire STAGE_31_OUT_1, STAGE_31_OUT_2;
       NOR2_X2 X_NOR_STAGE_31_1 (.A1(STAGE_30_OUT_1), .A2(STAGE_30_OUT_2), .ZN(STAGE_31_OUT_1));
       NOR2_X2 X_NOR_STAGE_31_2 (.A1(STAGE_30_OUT_1), .A2(STAGE_30_OUT_2), .ZN(STAGE_31_OUT_2));

       wire STAGE_32_OUT_1, STAGE_32_OUT_2;
       NOR2_X2 X_NOR_STAGE_32_1 (.A1(STAGE_31_OUT_1), .A2(STAGE_31_OUT_2), .ZN(STAGE_32_OUT_1));
       NOR2_X2 X_NOR_STAGE_32_2 (.A1(STAGE_31_OUT_1), .A2(STAGE_31_OUT_2), .ZN(STAGE_32_OUT_2));

       wire STAGE_33_OUT_1, STAGE_33_OUT_2;
       NOR2_X2 X_NOR_STAGE_33_1 (.A1(STAGE_32_OUT_1), .A2(STAGE_32_OUT_2), .ZN(STAGE_33_OUT_1));
       NOR2_X2 X_NOR_STAGE_33_2 (.A1(STAGE_32_OUT_1), .A2(STAGE_32_OUT_2), .ZN(STAGE_33_OUT_2));

       wire STAGE_34_OUT_1, STAGE_34_OUT_2;
       NOR2_X2 X_NOR_STAGE_34_1 (.A1(STAGE_33_OUT_1), .A2(STAGE_33_OUT_2), .ZN(STAGE_34_OUT_1));
       NOR2_X2 X_NOR_STAGE_34_2 (.A1(STAGE_33_OUT_1), .A2(STAGE_33_OUT_2), .ZN(STAGE_34_OUT_2));

       wire STAGE_35_OUT_1, STAGE_35_OUT_2;
       NOR2_X2 X_NOR_STAGE_35_1 (.A1(STAGE_34_OUT_1), .A2(STAGE_34_OUT_2), .ZN(STAGE_35_OUT_1));
       NOR2_X2 X_NOR_STAGE_35_2 (.A1(STAGE_34_OUT_1), .A2(STAGE_34_OUT_2), .ZN(STAGE_35_OUT_2));

       wire STAGE_36_OUT_1, STAGE_36_OUT_2;
       NOR2_X2 X_NOR_STAGE_36_1 (.A1(STAGE_35_OUT_1), .A2(STAGE_35_OUT_2), .ZN(STAGE_36_OUT_1));
       NOR2_X2 X_NOR_STAGE_36_2 (.A1(STAGE_35_OUT_1), .A2(STAGE_35_OUT_2), .ZN(STAGE_36_OUT_2));

       wire STAGE_37_OUT_1, STAGE_37_OUT_2;
       NOR2_X2 X_NOR_STAGE_37_1 (.A1(STAGE_36_OUT_1), .A2(STAGE_36_OUT_2), .ZN(STAGE_37_OUT_1));
       NOR2_X2 X_NOR_STAGE_37_2 (.A1(STAGE_36_OUT_1), .A2(STAGE_36_OUT_2), .ZN(STAGE_37_OUT_2));

       wire STAGE_38_OUT_1, STAGE_38_OUT_2;
       NOR2_X2 X_NOR_STAGE_38_1 (.A1(STAGE_37_OUT_1), .A2(STAGE_37_OUT_2), .ZN(STAGE_38_OUT_1));
       NOR2_X2 X_NOR_STAGE_38_2 (.A1(STAGE_37_OUT_1), .A2(STAGE_37_OUT_2), .ZN(STAGE_38_OUT_2));

       wire STAGE_39_OUT_1, STAGE_39_OUT_2;
       NOR2_X2 X_NOR_STAGE_39_1 (.A1(STAGE_38_OUT_1), .A2(STAGE_38_OUT_2), .ZN(STAGE_39_OUT_1));
       NOR2_X2 X_NOR_STAGE_39_2 (.A1(STAGE_38_OUT_1), .A2(STAGE_38_OUT_2), .ZN(STAGE_39_OUT_2));

       wire STAGE_40_OUT_1, STAGE_40_OUT_2;
       NOR2_X2 X_NOR_STAGE_40_1 (.A1(STAGE_39_OUT_1), .A2(STAGE_39_OUT_2), .ZN(STAGE_40_OUT_1));
       NOR2_X2 X_NOR_STAGE_40_2 (.A1(STAGE_39_OUT_1), .A2(STAGE_39_OUT_2), .ZN(STAGE_40_OUT_2));

       wire STAGE_41_OUT_1, STAGE_41_OUT_2;
       NOR2_X2 X_NOR_STAGE_41_1 (.A1(STAGE_40_OUT_1), .A2(STAGE_40_OUT_2), .ZN(STAGE_41_OUT_1));
       NOR2_X2 X_NOR_STAGE_41_2 (.A1(STAGE_40_OUT_1), .A2(STAGE_40_OUT_2), .ZN(STAGE_41_OUT_2));

       wire STAGE_42_OUT_1, STAGE_42_OUT_2;
       NOR2_X2 X_NOR_STAGE_42_1 (.A1(STAGE_41_OUT_1), .A2(STAGE_41_OUT_2), .ZN(STAGE_42_OUT_1));
       NOR2_X2 X_NOR_STAGE_42_2 (.A1(STAGE_41_OUT_1), .A2(STAGE_41_OUT_2), .ZN(STAGE_42_OUT_2));

       wire STAGE_43_OUT_1, STAGE_43_OUT_2;
       NOR2_X2 X_NOR_STAGE_43_1 (.A1(STAGE_42_OUT_1), .A2(STAGE_42_OUT_2), .ZN(STAGE_43_OUT_1));
       NOR2_X2 X_NOR_STAGE_43_2 (.A1(STAGE_42_OUT_1), .A2(STAGE_42_OUT_2), .ZN(STAGE_43_OUT_2));

       wire STAGE_44_OUT_1, STAGE_44_OUT_2;
       NOR2_X2 X_NOR_STAGE_44_1 (.A1(STAGE_43_OUT_1), .A2(STAGE_43_OUT_2), .ZN(STAGE_44_OUT_1));
       NOR2_X2 X_NOR_STAGE_44_2 (.A1(STAGE_43_OUT_1), .A2(STAGE_43_OUT_2), .ZN(STAGE_44_OUT_2));

       wire STAGE_45_OUT_1, STAGE_45_OUT_2;
       NOR2_X2 X_NOR_STAGE_45_1 (.A1(STAGE_44_OUT_1), .A2(STAGE_44_OUT_2), .ZN(STAGE_45_OUT_1));
       NOR2_X2 X_NOR_STAGE_45_2 (.A1(STAGE_44_OUT_1), .A2(STAGE_44_OUT_2), .ZN(STAGE_45_OUT_2));

       wire STAGE_46_OUT_1, STAGE_46_OUT_2;
       NOR2_X2 X_NOR_STAGE_46_1 (.A1(STAGE_45_OUT_1), .A2(STAGE_45_OUT_2), .ZN(STAGE_46_OUT_1));
       NOR2_X2 X_NOR_STAGE_46_2 (.A1(STAGE_45_OUT_1), .A2(STAGE_45_OUT_2), .ZN(STAGE_46_OUT_2));

       wire STAGE_47_OUT_1, STAGE_47_OUT_2;
       NOR2_X2 X_NOR_STAGE_47_1 (.A1(STAGE_46_OUT_1), .A2(STAGE_46_OUT_2), .ZN(STAGE_47_OUT_1));
       NOR2_X2 X_NOR_STAGE_47_2 (.A1(STAGE_46_OUT_1), .A2(STAGE_46_OUT_2), .ZN(STAGE_47_OUT_2));

       wire STAGE_48_OUT_1, STAGE_48_OUT_2;
       NOR2_X2 X_NOR_STAGE_48_1 (.A1(STAGE_47_OUT_1), .A2(STAGE_47_OUT_2), .ZN(STAGE_48_OUT_1));
       NOR2_X2 X_NOR_STAGE_48_2 (.A1(STAGE_47_OUT_1), .A2(STAGE_47_OUT_2), .ZN(STAGE_48_OUT_2));

       wire STAGE_49_OUT_1, STAGE_49_OUT_2;
       NOR2_X2 X_NOR_STAGE_49_1 (.A1(STAGE_48_OUT_1), .A2(STAGE_48_OUT_2), .ZN(STAGE_49_OUT_1));
       NOR2_X2 X_NOR_STAGE_49_2 (.A1(STAGE_48_OUT_1), .A2(STAGE_48_OUT_2), .ZN(STAGE_49_OUT_2));

       wire STAGE_50_OUT_1, STAGE_50_OUT_2;
       NOR2_X2 X_NOR_STAGE_50_1 (.A1(STAGE_49_OUT_1), .A2(STAGE_49_OUT_2), .ZN(STAGE_50_OUT_1));
       NOR2_X2 X_NOR_STAGE_50_2 (.A1(STAGE_49_OUT_1), .A2(STAGE_49_OUT_2), .ZN(STAGE_50_OUT_2));

       wire STAGE_51_OUT_1, STAGE_51_OUT_2;
       NOR2_X2 X_NOR_STAGE_51_1 (.A1(STAGE_50_OUT_1), .A2(STAGE_50_OUT_2), .ZN(STAGE_51_OUT_1));
       NOR2_X2 X_NOR_STAGE_51_2 (.A1(STAGE_50_OUT_1), .A2(STAGE_50_OUT_2), .ZN(STAGE_51_OUT_2));

       wire STAGE_52_OUT_1, STAGE_52_OUT_2;
       NOR2_X2 X_NOR_STAGE_52_1 (.A1(STAGE_51_OUT_1), .A2(STAGE_51_OUT_2), .ZN(STAGE_52_OUT_1));
       NOR2_X2 X_NOR_STAGE_52_2 (.A1(STAGE_51_OUT_1), .A2(STAGE_51_OUT_2), .ZN(STAGE_52_OUT_2));

       wire STAGE_53_OUT_1, STAGE_53_OUT_2;
       NOR2_X2 X_NOR_STAGE_53_1 (.A1(STAGE_52_OUT_1), .A2(STAGE_52_OUT_2), .ZN(OUT_Z1));
       NOR2_X2 X_NOR_STAGE_53_2 (.A1(STAGE_52_OUT_1), .A2(STAGE_52_OUT_2), .ZN(OUT_Z2));

endmodule
* circuit: nor inv chain
simulator lang=spice

*.PARAM pw=<sed>pw<sed>as
.PARAM supp=0.8V slope=0.1fs
.PARAM t_init0=0.1ns t_init1=0.174ns
.PARAM baseVal=0V peakVal=0.8V tend=1.0ns


.LIB /home/s11777724/involution_tool_library_files/backend/spice/fet.inc CMG

* main circuit
.INCLUDE /home/s11777724/involution_tool_library_files/backend/spice/cell/NOR2_X1.sp

**** SPECTRE Back Annotation
.option spef='/home/s11777724/JS/idm_evaluation/parallel_NOR_chains_50_stages/place_and_route/parallel_NOR_chains_100_stages_renamed.spef'
****

.TEMP 25
.OPTION
+ INGOLD=2
+ PARHIER=LOCAL
*+ POST=CSDF
+ PROBE
+ BRIEF
+ ACCURATE
+ ABSVAR=0.0001
+ DVDT=2
+ RELTOL=1e-11
*+ DELMAX=100fs
+ dc_pivot_check=yes

* vdd
VDD VDD GND 0.8v

VIN IN_A GND PWL 0ns baseVal t_init0 baseVal 't_init0+slope' peakVal t_init1 peakVal 't_init1+slope' baseVal
VIN IN_B GND PWL 0ns baseVal t_init0 baseVal 't_init0+slope' peakVal t_init1 peakVal 't_init1+slope' baseVal

* circuit under test
X_NOR_STAGE_0_1 IN_A IN_B  STAGE_0_OUT_1 VDD VDD GND GND NOR2_X2
X_NOR_STAGE_0_2 IN_A IN_B  STAGE_0_OUT_2 VDD VDD GND GND NOR2_X2

X_NOR_STAGE_1_1 STAGE_0_OUT_1 STAGE_0_OUT_2  A1 VDD VDD GND GND NOR2_X2
X_NOR_STAGE_1_2 STAGE_0_OUT_1 STAGE_0_OUT_2  A2 VDD VDD GND GND NOR2_X2

X_NOR_STAGE_2_1 A1 A2  STAGE_2_OUT_1 VDD VDD GND GND NOR2_X2
X_NOR_STAGE_2_2 A1 A2  STAGE_2_OUT_2 VDD VDD GND GND NOR2_X2

X_NOR_STAGE_3_1 STAGE_2_OUT_1 STAGE_2_OUT_2  STAGE_3_OUT_1 VDD VDD GND GND NOR2_X2
X_NOR_STAGE_3_2 STAGE_2_OUT_1 STAGE_2_OUT_2  STAGE_3_OUT_2 VDD VDD GND GND NOR2_X2

X_NOR_STAGE_4_1 STAGE_3_OUT_1 STAGE_3_OUT_2  STAGE_4_OUT_1 VDD VDD GND GND NOR2_X2
X_NOR_STAGE_4_2 STAGE_3_OUT_1 STAGE_3_OUT_2  STAGE_4_OUT_2 VDD VDD GND GND NOR2_X2

X_NOR_STAGE_5_1 STAGE_4_OUT_1 STAGE_4_OUT_2  STAGE_5_OUT_1 VDD VDD GND GND NOR2_X2
X_NOR_STAGE_5_2 STAGE_4_OUT_1 STAGE_4_OUT_2  STAGE_5_OUT_2 VDD VDD GND GND NOR2_X2

X_NOR_STAGE_6_1 STAGE_5_OUT_1 STAGE_5_OUT_2  STAGE_6_OUT_1 VDD VDD GND GND NOR2_X2
X_NOR_STAGE_6_2 STAGE_5_OUT_1 STAGE_5_OUT_2  STAGE_6_OUT_2 VDD VDD GND GND NOR2_X2

X_NOR_STAGE_7_1 STAGE_6_OUT_1 STAGE_6_OUT_2  STAGE_7_OUT_1 VDD VDD GND GND NOR2_X2
X_NOR_STAGE_7_2 STAGE_6_OUT_1 STAGE_6_OUT_2  STAGE_7_OUT_2 VDD VDD GND GND NOR2_X2

X_NOR_STAGE_8_1 STAGE_7_OUT_1 STAGE_7_OUT_2  STAGE_8_OUT_1 VDD VDD GND GND NOR2_X2
X_NOR_STAGE_8_2 STAGE_7_OUT_1 STAGE_7_OUT_2  STAGE_8_OUT_2 VDD VDD GND GND NOR2_X2

X_NOR_STAGE_9_1 STAGE_8_OUT_1 STAGE_8_OUT_2  STAGE_9_OUT_1 VDD VDD GND GND NOR2_X2
X_NOR_STAGE_9_2 STAGE_8_OUT_1 STAGE_8_OUT_2  STAGE_9_OUT_2 VDD VDD GND GND NOR2_X2

X_NOR_STAGE_10_1 STAGE_9_OUT_1 STAGE_9_OUT_2  STAGE_10_OUT_1 VDD VDD GND GND NOR2_X2
X_NOR_STAGE_10_2 STAGE_9_OUT_1 STAGE_9_OUT_2  STAGE_10_OUT_2 VDD VDD GND GND NOR2_X2

X_NOR_STAGE_11_1 STAGE_10_OUT_1 STAGE_10_OUT_2  STAGE_11_OUT_1 VDD VDD GND GND NOR2_X2
X_NOR_STAGE_11_2 STAGE_10_OUT_1 STAGE_10_OUT_2  STAGE_11_OUT_2 VDD VDD GND GND NOR2_X2

X_NOR_STAGE_12_1 STAGE_11_OUT_1 STAGE_11_OUT_2  STAGE_12_OUT_1 VDD VDD GND GND NOR2_X2
X_NOR_STAGE_12_2 STAGE_11_OUT_1 STAGE_11_OUT_2  STAGE_12_OUT_2 VDD VDD GND GND NOR2_X2

X_NOR_STAGE_13_1 STAGE_12_OUT_1 STAGE_12_OUT_2  STAGE_13_OUT_1 VDD VDD GND GND NOR2_X2
X_NOR_STAGE_13_2 STAGE_12_OUT_1 STAGE_12_OUT_2  STAGE_13_OUT_2 VDD VDD GND GND NOR2_X2

X_NOR_STAGE_14_1 STAGE_13_OUT_1 STAGE_13_OUT_2  STAGE_14_OUT_1 VDD VDD GND GND NOR2_X2
X_NOR_STAGE_14_2 STAGE_13_OUT_1 STAGE_13_OUT_2  STAGE_14_OUT_2 VDD VDD GND GND NOR2_X2

X_NOR_STAGE_15_1 STAGE_14_OUT_1 STAGE_14_OUT_2  STAGE_15_OUT_1 VDD VDD GND GND NOR2_X2
X_NOR_STAGE_15_2 STAGE_14_OUT_1 STAGE_14_OUT_2  STAGE_15_OUT_2 VDD VDD GND GND NOR2_X2

X_NOR_STAGE_16_1 STAGE_15_OUT_1 STAGE_15_OUT_2  STAGE_16_OUT_1 VDD VDD GND GND NOR2_X2
X_NOR_STAGE_16_2 STAGE_15_OUT_1 STAGE_15_OUT_2  STAGE_16_OUT_2 VDD VDD GND GND NOR2_X2

X_NOR_STAGE_17_1 STAGE_16_OUT_1 STAGE_16_OUT_2  STAGE_17_OUT_1 VDD VDD GND GND NOR2_X2
X_NOR_STAGE_17_2 STAGE_16_OUT_1 STAGE_16_OUT_2  STAGE_17_OUT_2 VDD VDD GND GND NOR2_X2

X_NOR_STAGE_18_1 STAGE_17_OUT_1 STAGE_17_OUT_2  STAGE_18_OUT_1 VDD VDD GND GND NOR2_X2
X_NOR_STAGE_18_2 STAGE_17_OUT_1 STAGE_17_OUT_2  STAGE_18_OUT_2 VDD VDD GND GND NOR2_X2

X_NOR_STAGE_19_1 STAGE_18_OUT_1 STAGE_18_OUT_2  STAGE_19_OUT_1 VDD VDD GND GND NOR2_X2
X_NOR_STAGE_19_2 STAGE_18_OUT_1 STAGE_18_OUT_2  STAGE_19_OUT_2 VDD VDD GND GND NOR2_X2

X_NOR_STAGE_20_1 STAGE_19_OUT_1 STAGE_19_OUT_2  STAGE_20_OUT_1 VDD VDD GND GND NOR2_X2
X_NOR_STAGE_20_2 STAGE_19_OUT_1 STAGE_19_OUT_2  STAGE_20_OUT_2 VDD VDD GND GND NOR2_X2

X_NOR_STAGE_21_1 STAGE_20_OUT_1 STAGE_20_OUT_2  STAGE_21_OUT_1 VDD VDD GND GND NOR2_X2
X_NOR_STAGE_21_2 STAGE_20_OUT_1 STAGE_20_OUT_2  STAGE_21_OUT_2 VDD VDD GND GND NOR2_X2

X_NOR_STAGE_22_1 STAGE_21_OUT_1 STAGE_21_OUT_2  STAGE_22_OUT_1 VDD VDD GND GND NOR2_X2
X_NOR_STAGE_22_2 STAGE_21_OUT_1 STAGE_21_OUT_2  STAGE_22_OUT_2 VDD VDD GND GND NOR2_X2

X_NOR_STAGE_23_1 STAGE_22_OUT_1 STAGE_22_OUT_2  STAGE_23_OUT_1 VDD VDD GND GND NOR2_X2
X_NOR_STAGE_23_2 STAGE_22_OUT_1 STAGE_22_OUT_2  STAGE_23_OUT_2 VDD VDD GND GND NOR2_X2

X_NOR_STAGE_24_1 STAGE_23_OUT_1 STAGE_23_OUT_2  STAGE_24_OUT_1 VDD VDD GND GND NOR2_X2
X_NOR_STAGE_24_2 STAGE_23_OUT_1 STAGE_23_OUT_2  STAGE_24_OUT_2 VDD VDD GND GND NOR2_X2

X_NOR_STAGE_25_1 STAGE_24_OUT_1 STAGE_24_OUT_2  STAGE_25_OUT_1 VDD VDD GND GND NOR2_X2
X_NOR_STAGE_25_2 STAGE_24_OUT_1 STAGE_24_OUT_2  STAGE_25_OUT_2 VDD VDD GND GND NOR2_X2

X_NOR_STAGE_26_1 STAGE_25_OUT_1 STAGE_25_OUT_2  STAGE_26_OUT_1 VDD VDD GND GND NOR2_X2
X_NOR_STAGE_26_2 STAGE_25_OUT_1 STAGE_25_OUT_2  STAGE_26_OUT_2 VDD VDD GND GND NOR2_X2

X_NOR_STAGE_27_1 STAGE_26_OUT_1 STAGE_26_OUT_2  STAGE_27_OUT_1 VDD VDD GND GND NOR2_X2
X_NOR_STAGE_27_2 STAGE_26_OUT_1 STAGE_26_OUT_2  STAGE_27_OUT_2 VDD VDD GND GND NOR2_X2

X_NOR_STAGE_28_1 STAGE_27_OUT_1 STAGE_27_OUT_2  STAGE_28_OUT_1 VDD VDD GND GND NOR2_X2
X_NOR_STAGE_28_2 STAGE_27_OUT_1 STAGE_27_OUT_2  STAGE_28_OUT_2 VDD VDD GND GND NOR2_X2

X_NOR_STAGE_29_1 STAGE_28_OUT_1 STAGE_28_OUT_2  STAGE_29_OUT_1 VDD VDD GND GND NOR2_X2
X_NOR_STAGE_29_2 STAGE_28_OUT_1 STAGE_28_OUT_2  STAGE_29_OUT_2 VDD VDD GND GND NOR2_X2

X_NOR_STAGE_30_1 STAGE_29_OUT_1 STAGE_29_OUT_2  STAGE_30_OUT_1 VDD VDD GND GND NOR2_X2
X_NOR_STAGE_30_2 STAGE_29_OUT_1 STAGE_29_OUT_2  STAGE_30_OUT_2 VDD VDD GND GND NOR2_X2

X_NOR_STAGE_31_1 STAGE_30_OUT_1 STAGE_30_OUT_2  STAGE_31_OUT_1 VDD VDD GND GND NOR2_X2
X_NOR_STAGE_31_2 STAGE_30_OUT_1 STAGE_30_OUT_2  STAGE_31_OUT_2 VDD VDD GND GND NOR2_X2

X_NOR_STAGE_32_1 STAGE_31_OUT_1 STAGE_31_OUT_2  STAGE_32_OUT_1 VDD VDD GND GND NOR2_X2
X_NOR_STAGE_32_2 STAGE_31_OUT_1 STAGE_31_OUT_2  STAGE_32_OUT_2 VDD VDD GND GND NOR2_X2

X_NOR_STAGE_33_1 STAGE_32_OUT_1 STAGE_32_OUT_2  STAGE_33_OUT_1 VDD VDD GND GND NOR2_X2
X_NOR_STAGE_33_2 STAGE_32_OUT_1 STAGE_32_OUT_2  STAGE_33_OUT_2 VDD VDD GND GND NOR2_X2

X_NOR_STAGE_34_1 STAGE_33_OUT_1 STAGE_33_OUT_2  STAGE_34_OUT_1 VDD VDD GND GND NOR2_X2
X_NOR_STAGE_34_2 STAGE_33_OUT_1 STAGE_33_OUT_2  STAGE_34_OUT_2 VDD VDD GND GND NOR2_X2

X_NOR_STAGE_35_1 STAGE_34_OUT_1 STAGE_34_OUT_2  STAGE_35_OUT_1 VDD VDD GND GND NOR2_X2
X_NOR_STAGE_35_2 STAGE_34_OUT_1 STAGE_34_OUT_2  STAGE_35_OUT_2 VDD VDD GND GND NOR2_X2

X_NOR_STAGE_36_1 STAGE_35_OUT_1 STAGE_35_OUT_2  STAGE_36_OUT_1 VDD VDD GND GND NOR2_X2
X_NOR_STAGE_36_2 STAGE_35_OUT_1 STAGE_35_OUT_2  STAGE_36_OUT_2 VDD VDD GND GND NOR2_X2

X_NOR_STAGE_37_1 STAGE_36_OUT_1 STAGE_36_OUT_2  STAGE_37_OUT_1 VDD VDD GND GND NOR2_X2
X_NOR_STAGE_37_2 STAGE_36_OUT_1 STAGE_36_OUT_2  STAGE_37_OUT_2 VDD VDD GND GND NOR2_X2

X_NOR_STAGE_38_1 STAGE_37_OUT_1 STAGE_37_OUT_2  STAGE_38_OUT_1 VDD VDD GND GND NOR2_X2
X_NOR_STAGE_38_2 STAGE_37_OUT_1 STAGE_37_OUT_2  STAGE_38_OUT_2 VDD VDD GND GND NOR2_X2

X_NOR_STAGE_39_1 STAGE_38_OUT_1 STAGE_38_OUT_2  STAGE_39_OUT_1 VDD VDD GND GND NOR2_X2
X_NOR_STAGE_39_2 STAGE_38_OUT_1 STAGE_38_OUT_2  STAGE_39_OUT_2 VDD VDD GND GND NOR2_X2

X_NOR_STAGE_40_1 STAGE_39_OUT_1 STAGE_39_OUT_2  STAGE_40_OUT_1 VDD VDD GND GND NOR2_X2
X_NOR_STAGE_40_2 STAGE_39_OUT_1 STAGE_39_OUT_2  STAGE_40_OUT_2 VDD VDD GND GND NOR2_X2

X_NOR_STAGE_41_1 STAGE_40_OUT_1 STAGE_40_OUT_2  STAGE_41_OUT_1 VDD VDD GND GND NOR2_X2
X_NOR_STAGE_41_2 STAGE_40_OUT_1 STAGE_40_OUT_2  STAGE_41_OUT_2 VDD VDD GND GND NOR2_X2

X_NOR_STAGE_42_1 STAGE_41_OUT_1 STAGE_41_OUT_2  STAGE_42_OUT_1 VDD VDD GND GND NOR2_X2
X_NOR_STAGE_42_2 STAGE_41_OUT_1 STAGE_41_OUT_2  STAGE_42_OUT_2 VDD VDD GND GND NOR2_X2

X_NOR_STAGE_43_1 STAGE_42_OUT_1 STAGE_42_OUT_2  STAGE_43_OUT_1 VDD VDD GND GND NOR2_X2
X_NOR_STAGE_43_2 STAGE_42_OUT_1 STAGE_42_OUT_2  STAGE_43_OUT_2 VDD VDD GND GND NOR2_X2

X_NOR_STAGE_44_1 STAGE_43_OUT_1 STAGE_43_OUT_2  STAGE_44_OUT_1 VDD VDD GND GND NOR2_X2
X_NOR_STAGE_44_2 STAGE_43_OUT_1 STAGE_43_OUT_2  STAGE_44_OUT_2 VDD VDD GND GND NOR2_X2

X_NOR_STAGE_45_1 STAGE_44_OUT_1 STAGE_44_OUT_2  STAGE_45_OUT_1 VDD VDD GND GND NOR2_X2
X_NOR_STAGE_45_2 STAGE_44_OUT_1 STAGE_44_OUT_2  STAGE_45_OUT_2 VDD VDD GND GND NOR2_X2

X_NOR_STAGE_46_1 STAGE_45_OUT_1 STAGE_45_OUT_2  STAGE_46_OUT_1 VDD VDD GND GND NOR2_X2
X_NOR_STAGE_46_2 STAGE_45_OUT_1 STAGE_45_OUT_2  STAGE_46_OUT_2 VDD VDD GND GND NOR2_X2

X_NOR_STAGE_47_1 STAGE_46_OUT_1 STAGE_46_OUT_2  STAGE_47_OUT_1 VDD VDD GND GND NOR2_X2
X_NOR_STAGE_47_2 STAGE_46_OUT_1 STAGE_46_OUT_2  STAGE_47_OUT_2 VDD VDD GND GND NOR2_X2

X_NOR_STAGE_48_1 STAGE_47_OUT_1 STAGE_47_OUT_2  STAGE_48_OUT_1 VDD VDD GND GND NOR2_X2
X_NOR_STAGE_48_2 STAGE_47_OUT_1 STAGE_47_OUT_2  STAGE_48_OUT_2 VDD VDD GND GND NOR2_X2

X_NOR_STAGE_49_1 STAGE_48_OUT_1 STAGE_48_OUT_2  STAGE_49_OUT_1 VDD VDD GND GND NOR2_X2
X_NOR_STAGE_49_2 STAGE_48_OUT_1 STAGE_48_OUT_2  STAGE_49_OUT_2 VDD VDD GND GND NOR2_X2

X_NOR_STAGE_50_1 STAGE_49_OUT_1 STAGE_49_OUT_2  STAGE_50_OUT_1 VDD VDD GND GND NOR2_X2
X_NOR_STAGE_50_2 STAGE_49_OUT_1 STAGE_49_OUT_2  STAGE_50_OUT_2 VDD VDD GND GND NOR2_X2

X_NOR_STAGE_51_1 STAGE_50_OUT_1 STAGE_50_OUT_2  STAGE_51_OUT_1 VDD VDD GND GND NOR2_X2
X_NOR_STAGE_51_2 STAGE_50_OUT_1 STAGE_50_OUT_2  STAGE_51_OUT_2 VDD VDD GND GND NOR2_X2

X_NOR_STAGE_52_1 STAGE_51_OUT_1 STAGE_51_OUT_2  STAGE_52_OUT_1 VDD VDD GND GND NOR2_X2
X_NOR_STAGE_52_2 STAGE_51_OUT_1 STAGE_51_OUT_2  STAGE_52_OUT_2 VDD VDD GND GND NOR2_X2

X_NOR_STAGE_53_1 STAGE_52_OUT_1 STAGE_52_OUT_2  STAGE_53_OUT_1 VDD VDD GND GND NOR2_X2
X_NOR_STAGE_53_2 STAGE_52_OUT_1 STAGE_52_OUT_2  STAGE_53_OUT_2 VDD VDD GND GND NOR2_X2

X_NOR_STAGE_54_1 STAGE_53_OUT_1 STAGE_53_OUT_2  STAGE_54_OUT_1 VDD VDD GND GND NOR2_X2
X_NOR_STAGE_54_2 STAGE_53_OUT_1 STAGE_53_OUT_2  STAGE_54_OUT_2 VDD VDD GND GND NOR2_X2

X_NOR_STAGE_55_1 STAGE_54_OUT_1 STAGE_54_OUT_2  STAGE_55_OUT_1 VDD VDD GND GND NOR2_X2
X_NOR_STAGE_55_2 STAGE_54_OUT_1 STAGE_54_OUT_2  STAGE_55_OUT_2 VDD VDD GND GND NOR2_X2

X_NOR_STAGE_56_1 STAGE_55_OUT_1 STAGE_55_OUT_2  STAGE_56_OUT_1 VDD VDD GND GND NOR2_X2
X_NOR_STAGE_56_2 STAGE_55_OUT_1 STAGE_55_OUT_2  STAGE_56_OUT_2 VDD VDD GND GND NOR2_X2

X_NOR_STAGE_57_1 STAGE_56_OUT_1 STAGE_56_OUT_2  STAGE_57_OUT_1 VDD VDD GND GND NOR2_X2
X_NOR_STAGE_57_2 STAGE_56_OUT_1 STAGE_56_OUT_2  STAGE_57_OUT_2 VDD VDD GND GND NOR2_X2

X_NOR_STAGE_58_1 STAGE_57_OUT_1 STAGE_57_OUT_2  STAGE_58_OUT_1 VDD VDD GND GND NOR2_X2
X_NOR_STAGE_58_2 STAGE_57_OUT_1 STAGE_57_OUT_2  STAGE_58_OUT_2 VDD VDD GND GND NOR2_X2

X_NOR_STAGE_59_1 STAGE_58_OUT_1 STAGE_58_OUT_2  STAGE_59_OUT_1 VDD VDD GND GND NOR2_X2
X_NOR_STAGE_59_2 STAGE_58_OUT_1 STAGE_58_OUT_2  STAGE_59_OUT_2 VDD VDD GND GND NOR2_X2

X_NOR_STAGE_60_1 STAGE_59_OUT_1 STAGE_59_OUT_2  STAGE_60_OUT_1 VDD VDD GND GND NOR2_X2
X_NOR_STAGE_60_2 STAGE_59_OUT_1 STAGE_59_OUT_2  STAGE_60_OUT_2 VDD VDD GND GND NOR2_X2

X_NOR_STAGE_61_1 STAGE_60_OUT_1 STAGE_60_OUT_2  STAGE_61_OUT_1 VDD VDD GND GND NOR2_X2
X_NOR_STAGE_61_2 STAGE_60_OUT_1 STAGE_60_OUT_2  STAGE_61_OUT_2 VDD VDD GND GND NOR2_X2

X_NOR_STAGE_62_1 STAGE_61_OUT_1 STAGE_61_OUT_2  STAGE_62_OUT_1 VDD VDD GND GND NOR2_X2
X_NOR_STAGE_62_2 STAGE_61_OUT_1 STAGE_61_OUT_2  STAGE_62_OUT_2 VDD VDD GND GND NOR2_X2

X_NOR_STAGE_63_1 STAGE_62_OUT_1 STAGE_62_OUT_2  STAGE_63_OUT_1 VDD VDD GND GND NOR2_X2
X_NOR_STAGE_63_2 STAGE_62_OUT_1 STAGE_62_OUT_2  STAGE_63_OUT_2 VDD VDD GND GND NOR2_X2

X_NOR_STAGE_64_1 STAGE_63_OUT_1 STAGE_63_OUT_2  STAGE_64_OUT_1 VDD VDD GND GND NOR2_X2
X_NOR_STAGE_64_2 STAGE_63_OUT_1 STAGE_63_OUT_2  STAGE_64_OUT_2 VDD VDD GND GND NOR2_X2

X_NOR_STAGE_65_1 STAGE_64_OUT_1 STAGE_64_OUT_2  STAGE_65_OUT_1 VDD VDD GND GND NOR2_X2
X_NOR_STAGE_65_2 STAGE_64_OUT_1 STAGE_64_OUT_2  STAGE_65_OUT_2 VDD VDD GND GND NOR2_X2

X_NOR_STAGE_66_1 STAGE_65_OUT_1 STAGE_65_OUT_2  STAGE_66_OUT_1 VDD VDD GND GND NOR2_X2
X_NOR_STAGE_66_2 STAGE_65_OUT_1 STAGE_65_OUT_2  STAGE_66_OUT_2 VDD VDD GND GND NOR2_X2

X_NOR_STAGE_67_1 STAGE_66_OUT_1 STAGE_66_OUT_2  STAGE_67_OUT_1 VDD VDD GND GND NOR2_X2
X_NOR_STAGE_67_2 STAGE_66_OUT_1 STAGE_66_OUT_2  STAGE_67_OUT_2 VDD VDD GND GND NOR2_X2

X_NOR_STAGE_68_1 STAGE_67_OUT_1 STAGE_67_OUT_2  STAGE_68_OUT_1 VDD VDD GND GND NOR2_X2
X_NOR_STAGE_68_2 STAGE_67_OUT_1 STAGE_67_OUT_2  STAGE_68_OUT_2 VDD VDD GND GND NOR2_X2

X_NOR_STAGE_69_1 STAGE_68_OUT_1 STAGE_68_OUT_2  STAGE_69_OUT_1 VDD VDD GND GND NOR2_X2
X_NOR_STAGE_69_2 STAGE_68_OUT_1 STAGE_68_OUT_2  STAGE_69_OUT_2 VDD VDD GND GND NOR2_X2

X_NOR_STAGE_70_1 STAGE_69_OUT_1 STAGE_69_OUT_2  STAGE_70_OUT_1 VDD VDD GND GND NOR2_X2
X_NOR_STAGE_70_2 STAGE_69_OUT_1 STAGE_69_OUT_2  STAGE_70_OUT_2 VDD VDD GND GND NOR2_X2

X_NOR_STAGE_71_1 STAGE_70_OUT_1 STAGE_70_OUT_2  STAGE_71_OUT_1 VDD VDD GND GND NOR2_X2
X_NOR_STAGE_71_2 STAGE_70_OUT_1 STAGE_70_OUT_2  STAGE_71_OUT_2 VDD VDD GND GND NOR2_X2

X_NOR_STAGE_72_1 STAGE_71_OUT_1 STAGE_71_OUT_2  STAGE_72_OUT_1 VDD VDD GND GND NOR2_X2
X_NOR_STAGE_72_2 STAGE_71_OUT_1 STAGE_71_OUT_2  STAGE_72_OUT_2 VDD VDD GND GND NOR2_X2

X_NOR_STAGE_73_1 STAGE_72_OUT_1 STAGE_72_OUT_2  STAGE_73_OUT_1 VDD VDD GND GND NOR2_X2
X_NOR_STAGE_73_2 STAGE_72_OUT_1 STAGE_72_OUT_2  STAGE_73_OUT_2 VDD VDD GND GND NOR2_X2

X_NOR_STAGE_74_1 STAGE_73_OUT_1 STAGE_73_OUT_2  STAGE_74_OUT_1 VDD VDD GND GND NOR2_X2
X_NOR_STAGE_74_2 STAGE_73_OUT_1 STAGE_73_OUT_2  STAGE_74_OUT_2 VDD VDD GND GND NOR2_X2

X_NOR_STAGE_75_1 STAGE_74_OUT_1 STAGE_74_OUT_2  STAGE_75_OUT_1 VDD VDD GND GND NOR2_X2
X_NOR_STAGE_75_2 STAGE_74_OUT_1 STAGE_74_OUT_2  STAGE_75_OUT_2 VDD VDD GND GND NOR2_X2

X_NOR_STAGE_76_1 STAGE_75_OUT_1 STAGE_75_OUT_2  STAGE_76_OUT_1 VDD VDD GND GND NOR2_X2
X_NOR_STAGE_76_2 STAGE_75_OUT_1 STAGE_75_OUT_2  STAGE_76_OUT_2 VDD VDD GND GND NOR2_X2

X_NOR_STAGE_77_1 STAGE_76_OUT_1 STAGE_76_OUT_2  STAGE_77_OUT_1 VDD VDD GND GND NOR2_X2
X_NOR_STAGE_77_2 STAGE_76_OUT_1 STAGE_76_OUT_2  STAGE_77_OUT_2 VDD VDD GND GND NOR2_X2

X_NOR_STAGE_78_1 STAGE_77_OUT_1 STAGE_77_OUT_2  STAGE_78_OUT_1 VDD VDD GND GND NOR2_X2
X_NOR_STAGE_78_2 STAGE_77_OUT_1 STAGE_77_OUT_2  STAGE_78_OUT_2 VDD VDD GND GND NOR2_X2

X_NOR_STAGE_79_1 STAGE_78_OUT_1 STAGE_78_OUT_2  STAGE_79_OUT_1 VDD VDD GND GND NOR2_X2
X_NOR_STAGE_79_2 STAGE_78_OUT_1 STAGE_78_OUT_2  STAGE_79_OUT_2 VDD VDD GND GND NOR2_X2

X_NOR_STAGE_80_1 STAGE_79_OUT_1 STAGE_79_OUT_2  STAGE_80_OUT_1 VDD VDD GND GND NOR2_X2
X_NOR_STAGE_80_2 STAGE_79_OUT_1 STAGE_79_OUT_2  STAGE_80_OUT_2 VDD VDD GND GND NOR2_X2

X_NOR_STAGE_81_1 STAGE_80_OUT_1 STAGE_80_OUT_2  STAGE_81_OUT_1 VDD VDD GND GND NOR2_X2
X_NOR_STAGE_81_2 STAGE_80_OUT_1 STAGE_80_OUT_2  STAGE_81_OUT_2 VDD VDD GND GND NOR2_X2

X_NOR_STAGE_82_1 STAGE_81_OUT_1 STAGE_81_OUT_2  STAGE_82_OUT_1 VDD VDD GND GND NOR2_X2
X_NOR_STAGE_82_2 STAGE_81_OUT_1 STAGE_81_OUT_2  STAGE_82_OUT_2 VDD VDD GND GND NOR2_X2

X_NOR_STAGE_83_1 STAGE_82_OUT_1 STAGE_82_OUT_2  STAGE_83_OUT_1 VDD VDD GND GND NOR2_X2
X_NOR_STAGE_83_2 STAGE_82_OUT_1 STAGE_82_OUT_2  STAGE_83_OUT_2 VDD VDD GND GND NOR2_X2

X_NOR_STAGE_84_1 STAGE_83_OUT_1 STAGE_83_OUT_2  STAGE_84_OUT_1 VDD VDD GND GND NOR2_X2
X_NOR_STAGE_84_2 STAGE_83_OUT_1 STAGE_83_OUT_2  STAGE_84_OUT_2 VDD VDD GND GND NOR2_X2

X_NOR_STAGE_85_1 STAGE_84_OUT_1 STAGE_84_OUT_2  STAGE_85_OUT_1 VDD VDD GND GND NOR2_X2
X_NOR_STAGE_85_2 STAGE_84_OUT_1 STAGE_84_OUT_2  STAGE_85_OUT_2 VDD VDD GND GND NOR2_X2

X_NOR_STAGE_86_1 STAGE_85_OUT_1 STAGE_85_OUT_2  STAGE_86_OUT_1 VDD VDD GND GND NOR2_X2
X_NOR_STAGE_86_2 STAGE_85_OUT_1 STAGE_85_OUT_2  STAGE_86_OUT_2 VDD VDD GND GND NOR2_X2

X_NOR_STAGE_87_1 STAGE_86_OUT_1 STAGE_86_OUT_2  STAGE_87_OUT_1 VDD VDD GND GND NOR2_X2
X_NOR_STAGE_87_2 STAGE_86_OUT_1 STAGE_86_OUT_2  STAGE_87_OUT_2 VDD VDD GND GND NOR2_X2

X_NOR_STAGE_88_1 STAGE_87_OUT_1 STAGE_87_OUT_2  STAGE_88_OUT_1 VDD VDD GND GND NOR2_X2
X_NOR_STAGE_88_2 STAGE_87_OUT_1 STAGE_87_OUT_2  STAGE_88_OUT_2 VDD VDD GND GND NOR2_X2

X_NOR_STAGE_89_1 STAGE_88_OUT_1 STAGE_88_OUT_2  STAGE_89_OUT_1 VDD VDD GND GND NOR2_X2
X_NOR_STAGE_89_2 STAGE_88_OUT_1 STAGE_88_OUT_2  STAGE_89_OUT_2 VDD VDD GND GND NOR2_X2

X_NOR_STAGE_90_1 STAGE_89_OUT_1 STAGE_89_OUT_2  STAGE_90_OUT_1 VDD VDD GND GND NOR2_X2
X_NOR_STAGE_90_2 STAGE_89_OUT_1 STAGE_89_OUT_2  STAGE_90_OUT_2 VDD VDD GND GND NOR2_X2

X_NOR_STAGE_91_1 STAGE_90_OUT_1 STAGE_90_OUT_2  STAGE_91_OUT_1 VDD VDD GND GND NOR2_X2
X_NOR_STAGE_91_2 STAGE_90_OUT_1 STAGE_90_OUT_2  STAGE_91_OUT_2 VDD VDD GND GND NOR2_X2

X_NOR_STAGE_92_1 STAGE_91_OUT_1 STAGE_91_OUT_2  STAGE_92_OUT_1 VDD VDD GND GND NOR2_X2
X_NOR_STAGE_92_2 STAGE_91_OUT_1 STAGE_91_OUT_2  STAGE_92_OUT_2 VDD VDD GND GND NOR2_X2

X_NOR_STAGE_93_1 STAGE_92_OUT_1 STAGE_92_OUT_2  STAGE_93_OUT_1 VDD VDD GND GND NOR2_X2
X_NOR_STAGE_93_2 STAGE_92_OUT_1 STAGE_92_OUT_2  STAGE_93_OUT_2 VDD VDD GND GND NOR2_X2

X_NOR_STAGE_94_1 STAGE_93_OUT_1 STAGE_93_OUT_2  STAGE_94_OUT_1 VDD VDD GND GND NOR2_X2
X_NOR_STAGE_94_2 STAGE_93_OUT_1 STAGE_93_OUT_2  STAGE_94_OUT_2 VDD VDD GND GND NOR2_X2

X_NOR_STAGE_95_1 STAGE_94_OUT_1 STAGE_94_OUT_2  STAGE_95_OUT_1 VDD VDD GND GND NOR2_X2
X_NOR_STAGE_95_2 STAGE_94_OUT_1 STAGE_94_OUT_2  STAGE_95_OUT_2 VDD VDD GND GND NOR2_X2

X_NOR_STAGE_96_1 STAGE_95_OUT_1 STAGE_95_OUT_2  STAGE_96_OUT_1 VDD VDD GND GND NOR2_X2
X_NOR_STAGE_96_2 STAGE_95_OUT_1 STAGE_95_OUT_2  STAGE_96_OUT_2 VDD VDD GND GND NOR2_X2

X_NOR_STAGE_97_1 STAGE_96_OUT_1 STAGE_96_OUT_2  STAGE_97_OUT_1 VDD VDD GND GND NOR2_X2
X_NOR_STAGE_97_2 STAGE_96_OUT_1 STAGE_96_OUT_2  STAGE_97_OUT_2 VDD VDD GND GND NOR2_X2

X_NOR_STAGE_98_1 STAGE_97_OUT_1 STAGE_97_OUT_2  STAGE_98_OUT_1 VDD VDD GND GND NOR2_X2
X_NOR_STAGE_98_2 STAGE_97_OUT_1 STAGE_97_OUT_2  STAGE_98_OUT_2 VDD VDD GND GND NOR2_X2

X_NOR_STAGE_99_1 STAGE_98_OUT_1 STAGE_98_OUT_2  STAGE_99_OUT_1 VDD VDD GND GND NOR2_X2
X_NOR_STAGE_99_2 STAGE_98_OUT_1 STAGE_98_OUT_2  STAGE_99_OUT_2 VDD VDD GND GND NOR2_X2

X_NOR_STAGE_100_1 STAGE_99_OUT_1 STAGE_99_OUT_2  STAGE_100_OUT_1 VDD VDD GND GND NOR2_X2
X_NOR_STAGE_100_2 STAGE_99_OUT_1 STAGE_99_OUT_2  STAGE_100_OUT_2 VDD VDD GND GND NOR2_X2

X_NOR_STAGE_101_1 STAGE_100_OUT_1 STAGE_100_OUT_2  Z1 VDD VDD GND GND NOR2_X2
X_NOR_STAGE_101_2 STAGE_100_OUT_1 STAGE_100_OUT_2  Z2 VDD VDD GND GND NOR2_X2

X_NOR_STAGE_102_1 Z1 Z2  STAGE_102_OUT_1 VDD VDD GND GND NOR2_X2
X_NOR_STAGE_102_2 Z1 Z2  STAGE_102_OUT_2 VDD VDD GND GND NOR2_X2

X_NOR_STAGE_103_1 STAGE_102_OUT_1 STAGE_102_OUT_2  STAGE_103_OUT_1 VDD VDD GND GND NOR2_X2
X_NOR_STAGE_103_2 STAGE_102_OUT_1 STAGE_102_OUT_2  STAGE_103_OUT_2 VDD VDD GND GND NOR2_X2

C_STAGE_103_TERM_1 STAGE_103_OUT_1 GND 0.01PF
C_STAGE_103_TERM_2 STAGE_103_OUT_2 GND 0.01PF


.PROBE TRAN V(A1) V(A2) V(Z1) V(Z2)
.TRAN 0.1ps tend
.END

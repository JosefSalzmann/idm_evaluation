* circuit: cgate_test
simulator lang=spice

*.PARAM pw=<sed>pw<sed>as
.PARAM supp=0.8V slope=0.1fs
.PARAM t_init0=0.1ns t_init1=0.174ns
.PARAM baseVal=0V peakVal=0.8V tend=8100.0ns


.LIB /home/s11777724/involution_tool_library_files/backend/spice/fet.inc CMG

* main circuit
.INCLUDE /home/s11777724/involution_tool_library_files/backend/spice/cell/BUF_X8.sp
.INCLUDE cgate.sp

**** SPECTRE Back Annotation
.option spef='/home/s11777724/JS/idm_evaluation/cgate_test/place_and_route/cgate_test_restitch.spef'
****

.TEMP 25
.OPTION
+ INGOLD=2
+ PARHIER=LOCAL
*+ POST=CSDF
+ PROBE
+ BRIEF
+ ACCURATE
+ ABSVAR=0.0001
+ DVDT=2
+ RELTOL=1e-11
*+ DELMAX=100fs
+ dc_pivot_check=yes

* vdd
VDD VDD GND 0.8v

.PARAM t_a_0=10ns
.PARAM t_a_1=20.0ns
.PARAM t_a_2=30ns
.PARAM t_a_3=40.0ns
.PARAM t_a_4=50ns
.PARAM t_a_5=60.0ns
.PARAM t_a_6=70ns
.PARAM t_a_7=80.0ns
.PARAM t_a_8=90ns
.PARAM t_a_9=100.0ns
.PARAM t_a_10=110ns
.PARAM t_a_11=120.0ns
.PARAM t_a_12=130ns
.PARAM t_a_13=140.0ns
.PARAM t_a_14=150ns
.PARAM t_a_15=160.0ns
.PARAM t_a_16=170ns
.PARAM t_a_17=180.0ns
.PARAM t_a_18=190ns
.PARAM t_a_19=200.0ns
.PARAM t_a_20=210ns
.PARAM t_a_21=220.0ns
.PARAM t_a_22=230ns
.PARAM t_a_23=240.0ns
.PARAM t_a_24=250ns
.PARAM t_a_25=260.0ns
.PARAM t_a_26=270ns
.PARAM t_a_27=280.0ns
.PARAM t_a_28=290ns
.PARAM t_a_29=300.0ns
.PARAM t_a_30=310ns
.PARAM t_a_31=320.0ns
.PARAM t_a_32=330ns
.PARAM t_a_33=340.0ns
.PARAM t_a_34=350ns
.PARAM t_a_35=360.0ns
.PARAM t_a_36=370ns
.PARAM t_a_37=380.0ns
.PARAM t_a_38=390ns
.PARAM t_a_39=400.0ns
.PARAM t_a_40=410ns
.PARAM t_a_41=420.0ns
.PARAM t_a_42=430ns
.PARAM t_a_43=440.0ns
.PARAM t_a_44=450ns
.PARAM t_a_45=460.0ns
.PARAM t_a_46=470ns
.PARAM t_a_47=480.0ns
.PARAM t_a_48=490ns
.PARAM t_a_49=500.0ns
.PARAM t_a_50=510ns
.PARAM t_a_51=520.0ns
.PARAM t_a_52=530ns
.PARAM t_a_53=540.0ns
.PARAM t_a_54=550ns
.PARAM t_a_55=560.0ns
.PARAM t_a_56=570ns
.PARAM t_a_57=580.0ns
.PARAM t_a_58=590ns
.PARAM t_a_59=600.0ns
.PARAM t_a_60=610ns
.PARAM t_a_61=620.0ns
.PARAM t_a_62=630ns
.PARAM t_a_63=640.0ns
.PARAM t_a_64=650ns
.PARAM t_a_65=660.0ns
.PARAM t_a_66=670ns
.PARAM t_a_67=680.0ns
.PARAM t_a_68=690ns
.PARAM t_a_69=700.0ns
.PARAM t_a_70=710ns
.PARAM t_a_71=720.0ns
.PARAM t_a_72=730ns
.PARAM t_a_73=740.0ns
.PARAM t_a_74=750ns
.PARAM t_a_75=760.0ns
.PARAM t_a_76=770ns
.PARAM t_a_77=780.0ns
.PARAM t_a_78=790ns
.PARAM t_a_79=800.0ns
.PARAM t_a_80=810ns
.PARAM t_a_81=820.0ns
.PARAM t_a_82=830ns
.PARAM t_a_83=840.0ns
.PARAM t_a_84=850ns
.PARAM t_a_85=860.0ns
.PARAM t_a_86=870ns
.PARAM t_a_87=880.0ns
.PARAM t_a_88=890ns
.PARAM t_a_89=900.0ns
.PARAM t_a_90=910ns
.PARAM t_a_91=920.0ns
.PARAM t_a_92=930ns
.PARAM t_a_93=940.0ns
.PARAM t_a_94=950ns
.PARAM t_a_95=960.0ns
.PARAM t_a_96=970ns
.PARAM t_a_97=980.0ns
.PARAM t_a_98=990ns
.PARAM t_a_99=1000.0ns
.PARAM t_a_100=1010ns
.PARAM t_a_101=1020.0ns
.PARAM t_a_102=1030ns
.PARAM t_a_103=1040.0ns
.PARAM t_a_104=1050ns
.PARAM t_a_105=1060.0ns
.PARAM t_a_106=1070ns
.PARAM t_a_107=1080.0ns
.PARAM t_a_108=1090ns
.PARAM t_a_109=1100.0ns
.PARAM t_a_110=1110ns
.PARAM t_a_111=1120.0ns
.PARAM t_a_112=1130ns
.PARAM t_a_113=1140.0ns
.PARAM t_a_114=1150ns
.PARAM t_a_115=1160.0ns
.PARAM t_a_116=1170ns
.PARAM t_a_117=1180.0ns
.PARAM t_a_118=1190ns
.PARAM t_a_119=1200.0ns
.PARAM t_a_120=1210ns
.PARAM t_a_121=1220.0ns
.PARAM t_a_122=1230ns
.PARAM t_a_123=1240.0ns
.PARAM t_a_124=1250ns
.PARAM t_a_125=1260.0ns
.PARAM t_a_126=1270ns
.PARAM t_a_127=1280.0ns
.PARAM t_a_128=1290ns
.PARAM t_a_129=1300.0ns
.PARAM t_a_130=1310ns
.PARAM t_a_131=1320.0ns
.PARAM t_a_132=1330ns
.PARAM t_a_133=1340.0ns
.PARAM t_a_134=1350ns
.PARAM t_a_135=1360.0ns
.PARAM t_a_136=1370ns
.PARAM t_a_137=1380.0ns
.PARAM t_a_138=1390ns
.PARAM t_a_139=1400.0ns
.PARAM t_a_140=1410ns
.PARAM t_a_141=1420.0ns
.PARAM t_a_142=1430ns
.PARAM t_a_143=1440.0ns
.PARAM t_a_144=1450ns
.PARAM t_a_145=1460.0ns
.PARAM t_a_146=1470ns
.PARAM t_a_147=1480.0ns
.PARAM t_a_148=1490ns
.PARAM t_a_149=1500.0ns
.PARAM t_a_150=1510ns
.PARAM t_a_151=1520.0ns
.PARAM t_a_152=1530ns
.PARAM t_a_153=1540.0ns
.PARAM t_a_154=1550ns
.PARAM t_a_155=1560.0ns
.PARAM t_a_156=1570ns
.PARAM t_a_157=1580.0ns
.PARAM t_a_158=1590ns
.PARAM t_a_159=1600.0ns
.PARAM t_a_160=1610ns
.PARAM t_a_161=1620.0ns
.PARAM t_a_162=1630ns
.PARAM t_a_163=1640.0ns
.PARAM t_a_164=1650ns
.PARAM t_a_165=1660.0ns
.PARAM t_a_166=1670ns
.PARAM t_a_167=1680.0ns
.PARAM t_a_168=1690ns
.PARAM t_a_169=1700.0ns
.PARAM t_a_170=1710ns
.PARAM t_a_171=1720.0ns
.PARAM t_a_172=1730ns
.PARAM t_a_173=1740.0ns
.PARAM t_a_174=1750ns
.PARAM t_a_175=1760.0ns
.PARAM t_a_176=1770ns
.PARAM t_a_177=1780.0ns
.PARAM t_a_178=1790ns
.PARAM t_a_179=1800.0ns
.PARAM t_a_180=1810ns
.PARAM t_a_181=1820.0ns
.PARAM t_a_182=1830ns
.PARAM t_a_183=1840.0ns
.PARAM t_a_184=1850ns
.PARAM t_a_185=1860.0ns
.PARAM t_a_186=1870ns
.PARAM t_a_187=1880.0ns
.PARAM t_a_188=1890ns
.PARAM t_a_189=1900.0ns
.PARAM t_a_190=1910ns
.PARAM t_a_191=1920.0ns
.PARAM t_a_192=1930ns
.PARAM t_a_193=1940.0ns
.PARAM t_a_194=1950ns
.PARAM t_a_195=1960.0ns
.PARAM t_a_196=1970ns
.PARAM t_a_197=1980.0ns
.PARAM t_a_198=1990ns
.PARAM t_a_199=2000.0ns
.PARAM t_a_200=2010ns
.PARAM t_a_201=2020.0ns
.PARAM t_a_202=2030ns
.PARAM t_a_203=2040.0ns
.PARAM t_a_204=2050ns
.PARAM t_a_205=2060.0ns
.PARAM t_a_206=2070ns
.PARAM t_a_207=2080.0ns
.PARAM t_a_208=2090ns
.PARAM t_a_209=2100.0ns
.PARAM t_a_210=2110ns
.PARAM t_a_211=2120.0ns
.PARAM t_a_212=2130ns
.PARAM t_a_213=2140.0ns
.PARAM t_a_214=2150ns
.PARAM t_a_215=2160.0ns
.PARAM t_a_216=2170ns
.PARAM t_a_217=2180.0ns
.PARAM t_a_218=2190ns
.PARAM t_a_219=2200.0ns
.PARAM t_a_220=2210ns
.PARAM t_a_221=2220.0ns
.PARAM t_a_222=2230ns
.PARAM t_a_223=2240.0ns
.PARAM t_a_224=2250ns
.PARAM t_a_225=2260.0ns
.PARAM t_a_226=2270ns
.PARAM t_a_227=2280.0ns
.PARAM t_a_228=2290ns
.PARAM t_a_229=2300.0ns
.PARAM t_a_230=2310ns
.PARAM t_a_231=2320.0ns
.PARAM t_a_232=2330ns
.PARAM t_a_233=2340.0ns
.PARAM t_a_234=2350ns
.PARAM t_a_235=2360.0ns
.PARAM t_a_236=2370ns
.PARAM t_a_237=2380.0ns
.PARAM t_a_238=2390ns
.PARAM t_a_239=2400.0ns
.PARAM t_a_240=2410ns
.PARAM t_a_241=2420.0ns
.PARAM t_a_242=2430ns
.PARAM t_a_243=2440.0ns
.PARAM t_a_244=2450ns
.PARAM t_a_245=2460.0ns
.PARAM t_a_246=2470ns
.PARAM t_a_247=2480.0ns
.PARAM t_a_248=2490ns
.PARAM t_a_249=2500.0ns
.PARAM t_a_250=2510ns
.PARAM t_a_251=2520.0ns
.PARAM t_a_252=2530ns
.PARAM t_a_253=2540.0ns
.PARAM t_a_254=2550ns
.PARAM t_a_255=2560.0ns
.PARAM t_a_256=2570ns
.PARAM t_a_257=2580.0ns
.PARAM t_a_258=2590ns
.PARAM t_a_259=2600.0ns
.PARAM t_a_260=2610ns
.PARAM t_a_261=2620.0ns
.PARAM t_a_262=2630ns
.PARAM t_a_263=2640.0ns
.PARAM t_a_264=2650ns
.PARAM t_a_265=2660.0ns
.PARAM t_a_266=2670ns
.PARAM t_a_267=2680.0ns
.PARAM t_a_268=2690ns
.PARAM t_a_269=2700.0ns
.PARAM t_a_270=2710ns
.PARAM t_a_271=2720.0ns
.PARAM t_a_272=2730ns
.PARAM t_a_273=2740.0ns
.PARAM t_a_274=2750ns
.PARAM t_a_275=2760.0ns
.PARAM t_a_276=2770ns
.PARAM t_a_277=2780.0ns
.PARAM t_a_278=2790ns
.PARAM t_a_279=2800.0ns
.PARAM t_a_280=2810ns
.PARAM t_a_281=2820.0ns
.PARAM t_a_282=2830ns
.PARAM t_a_283=2840.0ns
.PARAM t_a_284=2850ns
.PARAM t_a_285=2860.0ns
.PARAM t_a_286=2870ns
.PARAM t_a_287=2880.0ns
.PARAM t_a_288=2890ns
.PARAM t_a_289=2900.0ns
.PARAM t_a_290=2910ns
.PARAM t_a_291=2920.0ns
.PARAM t_a_292=2930ns
.PARAM t_a_293=2940.0ns
.PARAM t_a_294=2950ns
.PARAM t_a_295=2960.0ns
.PARAM t_a_296=2970ns
.PARAM t_a_297=2980.0ns
.PARAM t_a_298=2990ns
.PARAM t_a_299=3000.0ns
.PARAM t_a_300=3010ns
.PARAM t_a_301=3020.0ns
.PARAM t_a_302=3030ns
.PARAM t_a_303=3040.0ns
.PARAM t_a_304=3050ns
.PARAM t_a_305=3060.0ns
.PARAM t_a_306=3070ns
.PARAM t_a_307=3080.0ns
.PARAM t_a_308=3090ns
.PARAM t_a_309=3100.0ns
.PARAM t_a_310=3110ns
.PARAM t_a_311=3120.0ns
.PARAM t_a_312=3130ns
.PARAM t_a_313=3140.0ns
.PARAM t_a_314=3150ns
.PARAM t_a_315=3160.0ns
.PARAM t_a_316=3170ns
.PARAM t_a_317=3180.0ns
.PARAM t_a_318=3190ns
.PARAM t_a_319=3200.0ns
.PARAM t_a_320=3210ns
.PARAM t_a_321=3220.0ns
.PARAM t_a_322=3230ns
.PARAM t_a_323=3240.0ns
.PARAM t_a_324=3250ns
.PARAM t_a_325=3260.0ns
.PARAM t_a_326=3270ns
.PARAM t_a_327=3280.0ns
.PARAM t_a_328=3290ns
.PARAM t_a_329=3300.0ns
.PARAM t_a_330=3310ns
.PARAM t_a_331=3320.0ns
.PARAM t_a_332=3330ns
.PARAM t_a_333=3340.0ns
.PARAM t_a_334=3350ns
.PARAM t_a_335=3360.0ns
.PARAM t_a_336=3370ns
.PARAM t_a_337=3380.0ns
.PARAM t_a_338=3390ns
.PARAM t_a_339=3400.0ns
.PARAM t_a_340=3410ns
.PARAM t_a_341=3420.0ns
.PARAM t_a_342=3430ns
.PARAM t_a_343=3440.0ns
.PARAM t_a_344=3450ns
.PARAM t_a_345=3460.0ns
.PARAM t_a_346=3470ns
.PARAM t_a_347=3480.0ns
.PARAM t_a_348=3490ns
.PARAM t_a_349=3500.0ns
.PARAM t_a_350=3510ns
.PARAM t_a_351=3520.0ns
.PARAM t_a_352=3530ns
.PARAM t_a_353=3540.0ns
.PARAM t_a_354=3550ns
.PARAM t_a_355=3560.0ns
.PARAM t_a_356=3570ns
.PARAM t_a_357=3580.0ns
.PARAM t_a_358=3590ns
.PARAM t_a_359=3600.0ns
.PARAM t_a_360=3610ns
.PARAM t_a_361=3620.0ns
.PARAM t_a_362=3630ns
.PARAM t_a_363=3640.0ns
.PARAM t_a_364=3650ns
.PARAM t_a_365=3660.0ns
.PARAM t_a_366=3670ns
.PARAM t_a_367=3680.0ns
.PARAM t_a_368=3690ns
.PARAM t_a_369=3700.0ns
.PARAM t_a_370=3710ns
.PARAM t_a_371=3720.0ns
.PARAM t_a_372=3730ns
.PARAM t_a_373=3740.0ns
.PARAM t_a_374=3750ns
.PARAM t_a_375=3760.0ns
.PARAM t_a_376=3770ns
.PARAM t_a_377=3780.0ns
.PARAM t_a_378=3790ns
.PARAM t_a_379=3800.0ns
.PARAM t_a_380=3810ns
.PARAM t_a_381=3820.0ns
.PARAM t_a_382=3830ns
.PARAM t_a_383=3840.0ns
.PARAM t_a_384=3850ns
.PARAM t_a_385=3860.0ns
.PARAM t_a_386=3870ns
.PARAM t_a_387=3880.0ns
.PARAM t_a_388=3890ns
.PARAM t_a_389=3900.0ns
.PARAM t_a_390=3910ns
.PARAM t_a_391=3920.0ns
.PARAM t_a_392=3930ns
.PARAM t_a_393=3940.0ns
.PARAM t_a_394=3950ns
.PARAM t_a_395=3960.0ns
.PARAM t_a_396=3970ns
.PARAM t_a_397=3980.0ns
.PARAM t_a_398=3990ns
.PARAM t_a_399=4000.0ns
.PARAM t_a_400=4010ns
.PARAM t_a_401=4020.0ns
.PARAM t_a_402=4030ns
.PARAM t_a_403=4040.0ns
.PARAM t_a_404=4050ns
.PARAM t_a_405=4060.0ns
.PARAM t_a_406=4070ns
.PARAM t_a_407=4080.0ns
.PARAM t_a_408=4090ns
.PARAM t_a_409=4100.0ns
.PARAM t_a_410=4110ns
.PARAM t_a_411=4120.0ns
.PARAM t_a_412=4130ns
.PARAM t_a_413=4140.0ns
.PARAM t_a_414=4150ns
.PARAM t_a_415=4160.0ns
.PARAM t_a_416=4170ns
.PARAM t_a_417=4180.0ns
.PARAM t_a_418=4190ns
.PARAM t_a_419=4200.0ns
.PARAM t_a_420=4210ns
.PARAM t_a_421=4220.0ns
.PARAM t_a_422=4230ns
.PARAM t_a_423=4240.0ns
.PARAM t_a_424=4250ns
.PARAM t_a_425=4260.0ns
.PARAM t_a_426=4270ns
.PARAM t_a_427=4280.0ns
.PARAM t_a_428=4290ns
.PARAM t_a_429=4300.0ns
.PARAM t_a_430=4310ns
.PARAM t_a_431=4320.0ns
.PARAM t_a_432=4330ns
.PARAM t_a_433=4340.0ns
.PARAM t_a_434=4350ns
.PARAM t_a_435=4360.0ns
.PARAM t_a_436=4370ns
.PARAM t_a_437=4380.0ns
.PARAM t_a_438=4390ns
.PARAM t_a_439=4400.0ns
.PARAM t_a_440=4410ns
.PARAM t_a_441=4420.0ns
.PARAM t_a_442=4430ns
.PARAM t_a_443=4440.0ns
.PARAM t_a_444=4450ns
.PARAM t_a_445=4460.0ns
.PARAM t_a_446=4470ns
.PARAM t_a_447=4480.0ns
.PARAM t_a_448=4490ns
.PARAM t_a_449=4500.0ns
.PARAM t_a_450=4510ns
.PARAM t_a_451=4520.0ns
.PARAM t_a_452=4530ns
.PARAM t_a_453=4540.0ns
.PARAM t_a_454=4550ns
.PARAM t_a_455=4560.0ns
.PARAM t_a_456=4570ns
.PARAM t_a_457=4580.0ns
.PARAM t_a_458=4590ns
.PARAM t_a_459=4600.0ns
.PARAM t_a_460=4610ns
.PARAM t_a_461=4620.0ns
.PARAM t_a_462=4630ns
.PARAM t_a_463=4640.0ns
.PARAM t_a_464=4650ns
.PARAM t_a_465=4660.0ns
.PARAM t_a_466=4670ns
.PARAM t_a_467=4680.0ns
.PARAM t_a_468=4690ns
.PARAM t_a_469=4700.0ns
.PARAM t_a_470=4710ns
.PARAM t_a_471=4720.0ns
.PARAM t_a_472=4730ns
.PARAM t_a_473=4740.0ns
.PARAM t_a_474=4750ns
.PARAM t_a_475=4760.0ns
.PARAM t_a_476=4770ns
.PARAM t_a_477=4780.0ns
.PARAM t_a_478=4790ns
.PARAM t_a_479=4800.0ns
.PARAM t_a_480=4810ns
.PARAM t_a_481=4820.0ns
.PARAM t_a_482=4830ns
.PARAM t_a_483=4840.0ns
.PARAM t_a_484=4850ns
.PARAM t_a_485=4860.0ns
.PARAM t_a_486=4870ns
.PARAM t_a_487=4880.0ns
.PARAM t_a_488=4890ns
.PARAM t_a_489=4900.0ns
.PARAM t_a_490=4910ns
.PARAM t_a_491=4920.0ns
.PARAM t_a_492=4930ns
.PARAM t_a_493=4940.0ns
.PARAM t_a_494=4950ns
.PARAM t_a_495=4960.0ns
.PARAM t_a_496=4970ns
.PARAM t_a_497=4980.0ns
.PARAM t_a_498=4990ns
.PARAM t_a_499=5000.0ns
.PARAM t_a_500=5010ns
.PARAM t_a_501=5020.0ns
.PARAM t_a_502=5030ns
.PARAM t_a_503=5040.0ns
.PARAM t_a_504=5050ns
.PARAM t_a_505=5060.0ns
.PARAM t_a_506=5070ns
.PARAM t_a_507=5080.0ns
.PARAM t_a_508=5090ns
.PARAM t_a_509=5100.0ns
.PARAM t_a_510=5110ns
.PARAM t_a_511=5120.0ns
.PARAM t_a_512=5130ns
.PARAM t_a_513=5140.0ns
.PARAM t_a_514=5150ns
.PARAM t_a_515=5160.0ns
.PARAM t_a_516=5170ns
.PARAM t_a_517=5180.0ns
.PARAM t_a_518=5190ns
.PARAM t_a_519=5200.0ns
.PARAM t_a_520=5210ns
.PARAM t_a_521=5220.0ns
.PARAM t_a_522=5230ns
.PARAM t_a_523=5240.0ns
.PARAM t_a_524=5250ns
.PARAM t_a_525=5260.0ns
.PARAM t_a_526=5270ns
.PARAM t_a_527=5280.0ns
.PARAM t_a_528=5290ns
.PARAM t_a_529=5300.0ns
.PARAM t_a_530=5310ns
.PARAM t_a_531=5320.0ns
.PARAM t_a_532=5330ns
.PARAM t_a_533=5340.0ns
.PARAM t_a_534=5350ns
.PARAM t_a_535=5360.0ns
.PARAM t_a_536=5370ns
.PARAM t_a_537=5380.0ns
.PARAM t_a_538=5390ns
.PARAM t_a_539=5400.0ns
.PARAM t_a_540=5410ns
.PARAM t_a_541=5420.0ns
.PARAM t_a_542=5430ns
.PARAM t_a_543=5440.0ns
.PARAM t_a_544=5450ns
.PARAM t_a_545=5460.0ns
.PARAM t_a_546=5470ns
.PARAM t_a_547=5480.0ns
.PARAM t_a_548=5490ns
.PARAM t_a_549=5500.0ns
.PARAM t_a_550=5510ns
.PARAM t_a_551=5520.0ns
.PARAM t_a_552=5530ns
.PARAM t_a_553=5540.0ns
.PARAM t_a_554=5550ns
.PARAM t_a_555=5560.0ns
.PARAM t_a_556=5570ns
.PARAM t_a_557=5580.0ns
.PARAM t_a_558=5590ns
.PARAM t_a_559=5600.0ns
.PARAM t_a_560=5610ns
.PARAM t_a_561=5620.0ns
.PARAM t_a_562=5630ns
.PARAM t_a_563=5640.0ns
.PARAM t_a_564=5650ns
.PARAM t_a_565=5660.0ns
.PARAM t_a_566=5670ns
.PARAM t_a_567=5680.0ns
.PARAM t_a_568=5690ns
.PARAM t_a_569=5700.0ns
.PARAM t_a_570=5710ns
.PARAM t_a_571=5720.0ns
.PARAM t_a_572=5730ns
.PARAM t_a_573=5740.0ns
.PARAM t_a_574=5750ns
.PARAM t_a_575=5760.0ns
.PARAM t_a_576=5770ns
.PARAM t_a_577=5780.0ns
.PARAM t_a_578=5790ns
.PARAM t_a_579=5800.0ns
.PARAM t_a_580=5810ns
.PARAM t_a_581=5820.0ns
.PARAM t_a_582=5830ns
.PARAM t_a_583=5840.0ns
.PARAM t_a_584=5850ns
.PARAM t_a_585=5860.0ns
.PARAM t_a_586=5870ns
.PARAM t_a_587=5880.0ns
.PARAM t_a_588=5890ns
.PARAM t_a_589=5900.0ns
.PARAM t_a_590=5910ns
.PARAM t_a_591=5920.0ns
.PARAM t_a_592=5930ns
.PARAM t_a_593=5940.0ns
.PARAM t_a_594=5950ns
.PARAM t_a_595=5960.0ns
.PARAM t_a_596=5970ns
.PARAM t_a_597=5980.0ns
.PARAM t_a_598=5990ns
.PARAM t_a_599=6000.0ns
.PARAM t_a_600=6010ns
.PARAM t_a_601=6020.0ns
.PARAM t_a_602=6030ns
.PARAM t_a_603=6040.0ns
.PARAM t_a_604=6050ns
.PARAM t_a_605=6060.0ns
.PARAM t_a_606=6070ns
.PARAM t_a_607=6080.0ns
.PARAM t_a_608=6090ns
.PARAM t_a_609=6100.0ns
.PARAM t_a_610=6110ns
.PARAM t_a_611=6120.0ns
.PARAM t_a_612=6130ns
.PARAM t_a_613=6140.0ns
.PARAM t_a_614=6150ns
.PARAM t_a_615=6160.0ns
.PARAM t_a_616=6170ns
.PARAM t_a_617=6180.0ns
.PARAM t_a_618=6190ns
.PARAM t_a_619=6200.0ns
.PARAM t_a_620=6210ns
.PARAM t_a_621=6220.0ns
.PARAM t_a_622=6230ns
.PARAM t_a_623=6240.0ns
.PARAM t_a_624=6250ns
.PARAM t_a_625=6260.0ns
.PARAM t_a_626=6270ns
.PARAM t_a_627=6280.0ns
.PARAM t_a_628=6290ns
.PARAM t_a_629=6300.0ns
.PARAM t_a_630=6310ns
.PARAM t_a_631=6320.0ns
.PARAM t_a_632=6330ns
.PARAM t_a_633=6340.0ns
.PARAM t_a_634=6350ns
.PARAM t_a_635=6360.0ns
.PARAM t_a_636=6370ns
.PARAM t_a_637=6380.0ns
.PARAM t_a_638=6390ns
.PARAM t_a_639=6400.0ns
.PARAM t_a_640=6410ns
.PARAM t_a_641=6420.0ns
.PARAM t_a_642=6430ns
.PARAM t_a_643=6440.0ns
.PARAM t_a_644=6450ns
.PARAM t_a_645=6460.0ns
.PARAM t_a_646=6470ns
.PARAM t_a_647=6480.0ns
.PARAM t_a_648=6490ns
.PARAM t_a_649=6500.0ns
.PARAM t_a_650=6510ns
.PARAM t_a_651=6520.0ns
.PARAM t_a_652=6530ns
.PARAM t_a_653=6540.0ns
.PARAM t_a_654=6550ns
.PARAM t_a_655=6560.0ns
.PARAM t_a_656=6570ns
.PARAM t_a_657=6580.0ns
.PARAM t_a_658=6590ns
.PARAM t_a_659=6600.0ns
.PARAM t_a_660=6610ns
.PARAM t_a_661=6620.0ns
.PARAM t_a_662=6630ns
.PARAM t_a_663=6640.0ns
.PARAM t_a_664=6650ns
.PARAM t_a_665=6660.0ns
.PARAM t_a_666=6670ns
.PARAM t_a_667=6680.0ns
.PARAM t_a_668=6690ns
.PARAM t_a_669=6700.0ns
.PARAM t_a_670=6710ns
.PARAM t_a_671=6720.0ns
.PARAM t_a_672=6730ns
.PARAM t_a_673=6740.0ns
.PARAM t_a_674=6750ns
.PARAM t_a_675=6760.0ns
.PARAM t_a_676=6770ns
.PARAM t_a_677=6780.0ns
.PARAM t_a_678=6790ns
.PARAM t_a_679=6800.0ns
.PARAM t_a_680=6810ns
.PARAM t_a_681=6820.0ns
.PARAM t_a_682=6830ns
.PARAM t_a_683=6840.0ns
.PARAM t_a_684=6850ns
.PARAM t_a_685=6860.0ns
.PARAM t_a_686=6870ns
.PARAM t_a_687=6880.0ns
.PARAM t_a_688=6890ns
.PARAM t_a_689=6900.0ns
.PARAM t_a_690=6910ns
.PARAM t_a_691=6920.0ns
.PARAM t_a_692=6930ns
.PARAM t_a_693=6940.0ns
.PARAM t_a_694=6950ns
.PARAM t_a_695=6960.0ns
.PARAM t_a_696=6970ns
.PARAM t_a_697=6980.0ns
.PARAM t_a_698=6990ns
.PARAM t_a_699=7000.0ns
.PARAM t_a_700=7010ns
.PARAM t_a_701=7020.0ns
.PARAM t_a_702=7030ns
.PARAM t_a_703=7040.0ns
.PARAM t_a_704=7050ns
.PARAM t_a_705=7060.0ns
.PARAM t_a_706=7070ns
.PARAM t_a_707=7080.0ns
.PARAM t_a_708=7090ns
.PARAM t_a_709=7100.0ns
.PARAM t_a_710=7110ns
.PARAM t_a_711=7120.0ns
.PARAM t_a_712=7130ns
.PARAM t_a_713=7140.0ns
.PARAM t_a_714=7150ns
.PARAM t_a_715=7160.0ns
.PARAM t_a_716=7170ns
.PARAM t_a_717=7180.0ns
.PARAM t_a_718=7190ns
.PARAM t_a_719=7200.0ns
.PARAM t_a_720=7210ns
.PARAM t_a_721=7220.0ns
.PARAM t_a_722=7230ns
.PARAM t_a_723=7240.0ns
.PARAM t_a_724=7250ns
.PARAM t_a_725=7260.0ns
.PARAM t_a_726=7270ns
.PARAM t_a_727=7280.0ns
.PARAM t_a_728=7290ns
.PARAM t_a_729=7300.0ns
.PARAM t_a_730=7310ns
.PARAM t_a_731=7320.0ns
.PARAM t_a_732=7330ns
.PARAM t_a_733=7340.0ns
.PARAM t_a_734=7350ns
.PARAM t_a_735=7360.0ns
.PARAM t_a_736=7370ns
.PARAM t_a_737=7380.0ns
.PARAM t_a_738=7390ns
.PARAM t_a_739=7400.0ns
.PARAM t_a_740=7410ns
.PARAM t_a_741=7420.0ns
.PARAM t_a_742=7430ns
.PARAM t_a_743=7440.0ns
.PARAM t_a_744=7450ns
.PARAM t_a_745=7460.0ns
.PARAM t_a_746=7470ns
.PARAM t_a_747=7480.0ns
.PARAM t_a_748=7490ns
.PARAM t_a_749=7500.0ns
.PARAM t_a_750=7510ns
.PARAM t_a_751=7520.0ns
.PARAM t_a_752=7530ns
.PARAM t_a_753=7540.0ns
.PARAM t_a_754=7550ns
.PARAM t_a_755=7560.0ns
.PARAM t_a_756=7570ns
.PARAM t_a_757=7580.0ns
.PARAM t_a_758=7590ns
.PARAM t_a_759=7600.0ns
.PARAM t_a_760=7610ns
.PARAM t_a_761=7620.0ns
.PARAM t_a_762=7630ns
.PARAM t_a_763=7640.0ns
.PARAM t_a_764=7650ns
.PARAM t_a_765=7660.0ns
.PARAM t_a_766=7670ns
.PARAM t_a_767=7680.0ns
.PARAM t_a_768=7690ns
.PARAM t_a_769=7700.0ns
.PARAM t_a_770=7710ns
.PARAM t_a_771=7720.0ns
.PARAM t_a_772=7730ns
.PARAM t_a_773=7740.0ns
.PARAM t_a_774=7750ns
.PARAM t_a_775=7760.0ns
.PARAM t_a_776=7770ns
.PARAM t_a_777=7780.0ns
.PARAM t_a_778=7790ns
.PARAM t_a_779=7800.0ns
.PARAM t_a_780=7810ns
.PARAM t_a_781=7820.0ns
.PARAM t_a_782=7830ns
.PARAM t_a_783=7840.0ns
.PARAM t_a_784=7850ns
.PARAM t_a_785=7860.0ns
.PARAM t_a_786=7870ns
.PARAM t_a_787=7880.0ns
.PARAM t_a_788=7890ns
.PARAM t_a_789=7900.0ns
.PARAM t_a_790=7910ns
.PARAM t_a_791=7920.0ns
.PARAM t_a_792=7930ns
.PARAM t_a_793=7940.0ns
.PARAM t_a_794=7950ns
.PARAM t_a_795=7960.0ns
.PARAM t_a_796=7970ns
.PARAM t_a_797=7980.0ns
.PARAM t_a_798=7990ns
.PARAM t_a_799=8000.0ns
.PARAM t_b_0=9.9ns
.PARAM t_b_1=20.0ns
.PARAM t_b_2=29.9005ns
.PARAM t_b_3=40.0ns
.PARAM t_b_4=49.901ns
.PARAM t_b_5=60.0ns
.PARAM t_b_6=69.9015ns
.PARAM t_b_7=80.0ns
.PARAM t_b_8=89.902ns
.PARAM t_b_9=100.0ns
.PARAM t_b_10=109.9025ns
.PARAM t_b_11=120.0ns
.PARAM t_b_12=129.903ns
.PARAM t_b_13=140.0ns
.PARAM t_b_14=149.9035ns
.PARAM t_b_15=160.0ns
.PARAM t_b_16=169.904ns
.PARAM t_b_17=180.0ns
.PARAM t_b_18=189.9045ns
.PARAM t_b_19=200.0ns
.PARAM t_b_20=209.905ns
.PARAM t_b_21=220.0ns
.PARAM t_b_22=229.9055ns
.PARAM t_b_23=240.0ns
.PARAM t_b_24=249.906ns
.PARAM t_b_25=260.0ns
.PARAM t_b_26=269.9065ns
.PARAM t_b_27=280.0ns
.PARAM t_b_28=289.907ns
.PARAM t_b_29=300.0ns
.PARAM t_b_30=309.9075ns
.PARAM t_b_31=320.0ns
.PARAM t_b_32=329.908ns
.PARAM t_b_33=340.0ns
.PARAM t_b_34=349.9085ns
.PARAM t_b_35=360.0ns
.PARAM t_b_36=369.909ns
.PARAM t_b_37=380.0ns
.PARAM t_b_38=389.9095ns
.PARAM t_b_39=400.0ns
.PARAM t_b_40=409.91ns
.PARAM t_b_41=420.0ns
.PARAM t_b_42=429.9105ns
.PARAM t_b_43=440.0ns
.PARAM t_b_44=449.911ns
.PARAM t_b_45=460.0ns
.PARAM t_b_46=469.9115ns
.PARAM t_b_47=480.0ns
.PARAM t_b_48=489.912ns
.PARAM t_b_49=500.0ns
.PARAM t_b_50=509.9125ns
.PARAM t_b_51=520.0ns
.PARAM t_b_52=529.913ns
.PARAM t_b_53=540.0ns
.PARAM t_b_54=549.9135ns
.PARAM t_b_55=560.0ns
.PARAM t_b_56=569.914ns
.PARAM t_b_57=580.0ns
.PARAM t_b_58=589.9145ns
.PARAM t_b_59=600.0ns
.PARAM t_b_60=609.915ns
.PARAM t_b_61=620.0ns
.PARAM t_b_62=629.9155ns
.PARAM t_b_63=640.0ns
.PARAM t_b_64=649.916ns
.PARAM t_b_65=660.0ns
.PARAM t_b_66=669.9165ns
.PARAM t_b_67=680.0ns
.PARAM t_b_68=689.917ns
.PARAM t_b_69=700.0ns
.PARAM t_b_70=709.9175ns
.PARAM t_b_71=720.0ns
.PARAM t_b_72=729.918ns
.PARAM t_b_73=740.0ns
.PARAM t_b_74=749.9185ns
.PARAM t_b_75=760.0ns
.PARAM t_b_76=769.919ns
.PARAM t_b_77=780.0ns
.PARAM t_b_78=789.9195ns
.PARAM t_b_79=800.0ns
.PARAM t_b_80=809.92ns
.PARAM t_b_81=820.0ns
.PARAM t_b_82=829.9205ns
.PARAM t_b_83=840.0ns
.PARAM t_b_84=849.921ns
.PARAM t_b_85=860.0ns
.PARAM t_b_86=869.9215ns
.PARAM t_b_87=880.0ns
.PARAM t_b_88=889.922ns
.PARAM t_b_89=900.0ns
.PARAM t_b_90=909.9225ns
.PARAM t_b_91=920.0ns
.PARAM t_b_92=929.923ns
.PARAM t_b_93=940.0ns
.PARAM t_b_94=949.9235ns
.PARAM t_b_95=960.0ns
.PARAM t_b_96=969.924ns
.PARAM t_b_97=980.0ns
.PARAM t_b_98=989.9245ns
.PARAM t_b_99=1000.0ns
.PARAM t_b_100=1009.925ns
.PARAM t_b_101=1020.0ns
.PARAM t_b_102=1029.9255ns
.PARAM t_b_103=1040.0ns
.PARAM t_b_104=1049.926ns
.PARAM t_b_105=1060.0ns
.PARAM t_b_106=1069.9265ns
.PARAM t_b_107=1080.0ns
.PARAM t_b_108=1089.927ns
.PARAM t_b_109=1100.0ns
.PARAM t_b_110=1109.9275ns
.PARAM t_b_111=1120.0ns
.PARAM t_b_112=1129.928ns
.PARAM t_b_113=1140.0ns
.PARAM t_b_114=1149.9285ns
.PARAM t_b_115=1160.0ns
.PARAM t_b_116=1169.929ns
.PARAM t_b_117=1180.0ns
.PARAM t_b_118=1189.9295ns
.PARAM t_b_119=1200.0ns
.PARAM t_b_120=1209.93ns
.PARAM t_b_121=1220.0ns
.PARAM t_b_122=1229.9305ns
.PARAM t_b_123=1240.0ns
.PARAM t_b_124=1249.931ns
.PARAM t_b_125=1260.0ns
.PARAM t_b_126=1269.9315ns
.PARAM t_b_127=1280.0ns
.PARAM t_b_128=1289.932ns
.PARAM t_b_129=1300.0ns
.PARAM t_b_130=1309.9325ns
.PARAM t_b_131=1320.0ns
.PARAM t_b_132=1329.933ns
.PARAM t_b_133=1340.0ns
.PARAM t_b_134=1349.9335ns
.PARAM t_b_135=1360.0ns
.PARAM t_b_136=1369.934ns
.PARAM t_b_137=1380.0ns
.PARAM t_b_138=1389.9345ns
.PARAM t_b_139=1400.0ns
.PARAM t_b_140=1409.935ns
.PARAM t_b_141=1420.0ns
.PARAM t_b_142=1429.9355ns
.PARAM t_b_143=1440.0ns
.PARAM t_b_144=1449.936ns
.PARAM t_b_145=1460.0ns
.PARAM t_b_146=1469.9365ns
.PARAM t_b_147=1480.0ns
.PARAM t_b_148=1489.937ns
.PARAM t_b_149=1500.0ns
.PARAM t_b_150=1509.9375ns
.PARAM t_b_151=1520.0ns
.PARAM t_b_152=1529.938ns
.PARAM t_b_153=1540.0ns
.PARAM t_b_154=1549.9385ns
.PARAM t_b_155=1560.0ns
.PARAM t_b_156=1569.939ns
.PARAM t_b_157=1580.0ns
.PARAM t_b_158=1589.9395ns
.PARAM t_b_159=1600.0ns
.PARAM t_b_160=1609.94ns
.PARAM t_b_161=1620.0ns
.PARAM t_b_162=1629.9405ns
.PARAM t_b_163=1640.0ns
.PARAM t_b_164=1649.941ns
.PARAM t_b_165=1660.0ns
.PARAM t_b_166=1669.9415ns
.PARAM t_b_167=1680.0ns
.PARAM t_b_168=1689.942ns
.PARAM t_b_169=1700.0ns
.PARAM t_b_170=1709.9425ns
.PARAM t_b_171=1720.0ns
.PARAM t_b_172=1729.943ns
.PARAM t_b_173=1740.0ns
.PARAM t_b_174=1749.9435ns
.PARAM t_b_175=1760.0ns
.PARAM t_b_176=1769.944ns
.PARAM t_b_177=1780.0ns
.PARAM t_b_178=1789.9445ns
.PARAM t_b_179=1800.0ns
.PARAM t_b_180=1809.945ns
.PARAM t_b_181=1820.0ns
.PARAM t_b_182=1829.9455ns
.PARAM t_b_183=1840.0ns
.PARAM t_b_184=1849.946ns
.PARAM t_b_185=1860.0ns
.PARAM t_b_186=1869.9465ns
.PARAM t_b_187=1880.0ns
.PARAM t_b_188=1889.947ns
.PARAM t_b_189=1900.0ns
.PARAM t_b_190=1909.9475ns
.PARAM t_b_191=1920.0ns
.PARAM t_b_192=1929.948ns
.PARAM t_b_193=1940.0ns
.PARAM t_b_194=1949.9485ns
.PARAM t_b_195=1960.0ns
.PARAM t_b_196=1969.949ns
.PARAM t_b_197=1980.0ns
.PARAM t_b_198=1989.9495ns
.PARAM t_b_199=2000.0ns
.PARAM t_b_200=2009.95ns
.PARAM t_b_201=2020.0ns
.PARAM t_b_202=2029.9505ns
.PARAM t_b_203=2040.0ns
.PARAM t_b_204=2049.951ns
.PARAM t_b_205=2060.0ns
.PARAM t_b_206=2069.9515ns
.PARAM t_b_207=2080.0ns
.PARAM t_b_208=2089.952ns
.PARAM t_b_209=2100.0ns
.PARAM t_b_210=2109.9525ns
.PARAM t_b_211=2120.0ns
.PARAM t_b_212=2129.953ns
.PARAM t_b_213=2140.0ns
.PARAM t_b_214=2149.9535ns
.PARAM t_b_215=2160.0ns
.PARAM t_b_216=2169.954ns
.PARAM t_b_217=2180.0ns
.PARAM t_b_218=2189.9545ns
.PARAM t_b_219=2200.0ns
.PARAM t_b_220=2209.955ns
.PARAM t_b_221=2220.0ns
.PARAM t_b_222=2229.9555ns
.PARAM t_b_223=2240.0ns
.PARAM t_b_224=2249.956ns
.PARAM t_b_225=2260.0ns
.PARAM t_b_226=2269.9565ns
.PARAM t_b_227=2280.0ns
.PARAM t_b_228=2289.957ns
.PARAM t_b_229=2300.0ns
.PARAM t_b_230=2309.9575ns
.PARAM t_b_231=2320.0ns
.PARAM t_b_232=2329.958ns
.PARAM t_b_233=2340.0ns
.PARAM t_b_234=2349.9585ns
.PARAM t_b_235=2360.0ns
.PARAM t_b_236=2369.959ns
.PARAM t_b_237=2380.0ns
.PARAM t_b_238=2389.9595ns
.PARAM t_b_239=2400.0ns
.PARAM t_b_240=2409.96ns
.PARAM t_b_241=2420.0ns
.PARAM t_b_242=2429.9605ns
.PARAM t_b_243=2440.0ns
.PARAM t_b_244=2449.961ns
.PARAM t_b_245=2460.0ns
.PARAM t_b_246=2469.9615ns
.PARAM t_b_247=2480.0ns
.PARAM t_b_248=2489.962ns
.PARAM t_b_249=2500.0ns
.PARAM t_b_250=2509.9625ns
.PARAM t_b_251=2520.0ns
.PARAM t_b_252=2529.963ns
.PARAM t_b_253=2540.0ns
.PARAM t_b_254=2549.9635ns
.PARAM t_b_255=2560.0ns
.PARAM t_b_256=2569.964ns
.PARAM t_b_257=2580.0ns
.PARAM t_b_258=2589.9645ns
.PARAM t_b_259=2600.0ns
.PARAM t_b_260=2609.965ns
.PARAM t_b_261=2620.0ns
.PARAM t_b_262=2629.9655ns
.PARAM t_b_263=2640.0ns
.PARAM t_b_264=2649.966ns
.PARAM t_b_265=2660.0ns
.PARAM t_b_266=2669.9665ns
.PARAM t_b_267=2680.0ns
.PARAM t_b_268=2689.967ns
.PARAM t_b_269=2700.0ns
.PARAM t_b_270=2709.9675ns
.PARAM t_b_271=2720.0ns
.PARAM t_b_272=2729.968ns
.PARAM t_b_273=2740.0ns
.PARAM t_b_274=2749.9685ns
.PARAM t_b_275=2760.0ns
.PARAM t_b_276=2769.969ns
.PARAM t_b_277=2780.0ns
.PARAM t_b_278=2789.9695ns
.PARAM t_b_279=2800.0ns
.PARAM t_b_280=2809.97ns
.PARAM t_b_281=2820.0ns
.PARAM t_b_282=2829.9705ns
.PARAM t_b_283=2840.0ns
.PARAM t_b_284=2849.971ns
.PARAM t_b_285=2860.0ns
.PARAM t_b_286=2869.9715ns
.PARAM t_b_287=2880.0ns
.PARAM t_b_288=2889.972ns
.PARAM t_b_289=2900.0ns
.PARAM t_b_290=2909.9725ns
.PARAM t_b_291=2920.0ns
.PARAM t_b_292=2929.973ns
.PARAM t_b_293=2940.0ns
.PARAM t_b_294=2949.9735ns
.PARAM t_b_295=2960.0ns
.PARAM t_b_296=2969.974ns
.PARAM t_b_297=2980.0ns
.PARAM t_b_298=2989.9745ns
.PARAM t_b_299=3000.0ns
.PARAM t_b_300=3009.975ns
.PARAM t_b_301=3020.0ns
.PARAM t_b_302=3029.9755ns
.PARAM t_b_303=3040.0ns
.PARAM t_b_304=3049.976ns
.PARAM t_b_305=3060.0ns
.PARAM t_b_306=3069.9765ns
.PARAM t_b_307=3080.0ns
.PARAM t_b_308=3089.977ns
.PARAM t_b_309=3100.0ns
.PARAM t_b_310=3109.9775ns
.PARAM t_b_311=3120.0ns
.PARAM t_b_312=3129.978ns
.PARAM t_b_313=3140.0ns
.PARAM t_b_314=3149.9785ns
.PARAM t_b_315=3160.0ns
.PARAM t_b_316=3169.979ns
.PARAM t_b_317=3180.0ns
.PARAM t_b_318=3189.9795ns
.PARAM t_b_319=3200.0ns
.PARAM t_b_320=3209.98ns
.PARAM t_b_321=3220.0ns
.PARAM t_b_322=3229.9805ns
.PARAM t_b_323=3240.0ns
.PARAM t_b_324=3249.981ns
.PARAM t_b_325=3260.0ns
.PARAM t_b_326=3269.9815ns
.PARAM t_b_327=3280.0ns
.PARAM t_b_328=3289.982ns
.PARAM t_b_329=3300.0ns
.PARAM t_b_330=3309.9825ns
.PARAM t_b_331=3320.0ns
.PARAM t_b_332=3329.983ns
.PARAM t_b_333=3340.0ns
.PARAM t_b_334=3349.9835ns
.PARAM t_b_335=3360.0ns
.PARAM t_b_336=3369.984ns
.PARAM t_b_337=3380.0ns
.PARAM t_b_338=3389.9845ns
.PARAM t_b_339=3400.0ns
.PARAM t_b_340=3409.985ns
.PARAM t_b_341=3420.0ns
.PARAM t_b_342=3429.9855ns
.PARAM t_b_343=3440.0ns
.PARAM t_b_344=3449.986ns
.PARAM t_b_345=3460.0ns
.PARAM t_b_346=3469.9865ns
.PARAM t_b_347=3480.0ns
.PARAM t_b_348=3489.987ns
.PARAM t_b_349=3500.0ns
.PARAM t_b_350=3509.9875ns
.PARAM t_b_351=3520.0ns
.PARAM t_b_352=3529.988ns
.PARAM t_b_353=3540.0ns
.PARAM t_b_354=3549.9885ns
.PARAM t_b_355=3560.0ns
.PARAM t_b_356=3569.989ns
.PARAM t_b_357=3580.0ns
.PARAM t_b_358=3589.9895ns
.PARAM t_b_359=3600.0ns
.PARAM t_b_360=3609.99ns
.PARAM t_b_361=3620.0ns
.PARAM t_b_362=3629.9905ns
.PARAM t_b_363=3640.0ns
.PARAM t_b_364=3649.991ns
.PARAM t_b_365=3660.0ns
.PARAM t_b_366=3669.9915ns
.PARAM t_b_367=3680.0ns
.PARAM t_b_368=3689.992ns
.PARAM t_b_369=3700.0ns
.PARAM t_b_370=3709.9925ns
.PARAM t_b_371=3720.0ns
.PARAM t_b_372=3729.993ns
.PARAM t_b_373=3740.0ns
.PARAM t_b_374=3749.9935ns
.PARAM t_b_375=3760.0ns
.PARAM t_b_376=3769.994ns
.PARAM t_b_377=3780.0ns
.PARAM t_b_378=3789.9945ns
.PARAM t_b_379=3800.0ns
.PARAM t_b_380=3809.995ns
.PARAM t_b_381=3820.0ns
.PARAM t_b_382=3829.9955ns
.PARAM t_b_383=3840.0ns
.PARAM t_b_384=3849.996ns
.PARAM t_b_385=3860.0ns
.PARAM t_b_386=3869.9965ns
.PARAM t_b_387=3880.0ns
.PARAM t_b_388=3889.997ns
.PARAM t_b_389=3900.0ns
.PARAM t_b_390=3909.9975ns
.PARAM t_b_391=3920.0ns
.PARAM t_b_392=3929.998ns
.PARAM t_b_393=3940.0ns
.PARAM t_b_394=3949.9985ns
.PARAM t_b_395=3960.0ns
.PARAM t_b_396=3969.999ns
.PARAM t_b_397=3980.0ns
.PARAM t_b_398=3989.9995ns
.PARAM t_b_399=4000.0ns
.PARAM t_b_400=4010.0ns
.PARAM t_b_401=4020.0ns
.PARAM t_b_402=4030.0005ns
.PARAM t_b_403=4040.0ns
.PARAM t_b_404=4050.001ns
.PARAM t_b_405=4060.0ns
.PARAM t_b_406=4070.0015ns
.PARAM t_b_407=4080.0ns
.PARAM t_b_408=4090.002ns
.PARAM t_b_409=4100.0ns
.PARAM t_b_410=4110.0025ns
.PARAM t_b_411=4120.0ns
.PARAM t_b_412=4130.003ns
.PARAM t_b_413=4140.0ns
.PARAM t_b_414=4150.0035ns
.PARAM t_b_415=4160.0ns
.PARAM t_b_416=4170.004ns
.PARAM t_b_417=4180.0ns
.PARAM t_b_418=4190.0045ns
.PARAM t_b_419=4200.0ns
.PARAM t_b_420=4210.005ns
.PARAM t_b_421=4220.0ns
.PARAM t_b_422=4230.0055ns
.PARAM t_b_423=4240.0ns
.PARAM t_b_424=4250.006ns
.PARAM t_b_425=4260.0ns
.PARAM t_b_426=4270.0065ns
.PARAM t_b_427=4280.0ns
.PARAM t_b_428=4290.007ns
.PARAM t_b_429=4300.0ns
.PARAM t_b_430=4310.0075ns
.PARAM t_b_431=4320.0ns
.PARAM t_b_432=4330.008ns
.PARAM t_b_433=4340.0ns
.PARAM t_b_434=4350.0085ns
.PARAM t_b_435=4360.0ns
.PARAM t_b_436=4370.009ns
.PARAM t_b_437=4380.0ns
.PARAM t_b_438=4390.0095ns
.PARAM t_b_439=4400.0ns
.PARAM t_b_440=4410.01ns
.PARAM t_b_441=4420.0ns
.PARAM t_b_442=4430.0105ns
.PARAM t_b_443=4440.0ns
.PARAM t_b_444=4450.011ns
.PARAM t_b_445=4460.0ns
.PARAM t_b_446=4470.0115ns
.PARAM t_b_447=4480.0ns
.PARAM t_b_448=4490.012ns
.PARAM t_b_449=4500.0ns
.PARAM t_b_450=4510.0125ns
.PARAM t_b_451=4520.0ns
.PARAM t_b_452=4530.013ns
.PARAM t_b_453=4540.0ns
.PARAM t_b_454=4550.0135ns
.PARAM t_b_455=4560.0ns
.PARAM t_b_456=4570.014ns
.PARAM t_b_457=4580.0ns
.PARAM t_b_458=4590.0145ns
.PARAM t_b_459=4600.0ns
.PARAM t_b_460=4610.015ns
.PARAM t_b_461=4620.0ns
.PARAM t_b_462=4630.0155ns
.PARAM t_b_463=4640.0ns
.PARAM t_b_464=4650.016ns
.PARAM t_b_465=4660.0ns
.PARAM t_b_466=4670.0165ns
.PARAM t_b_467=4680.0ns
.PARAM t_b_468=4690.017ns
.PARAM t_b_469=4700.0ns
.PARAM t_b_470=4710.0175ns
.PARAM t_b_471=4720.0ns
.PARAM t_b_472=4730.018ns
.PARAM t_b_473=4740.0ns
.PARAM t_b_474=4750.0185ns
.PARAM t_b_475=4760.0ns
.PARAM t_b_476=4770.019ns
.PARAM t_b_477=4780.0ns
.PARAM t_b_478=4790.0195ns
.PARAM t_b_479=4800.0ns
.PARAM t_b_480=4810.02ns
.PARAM t_b_481=4820.0ns
.PARAM t_b_482=4830.0205ns
.PARAM t_b_483=4840.0ns
.PARAM t_b_484=4850.021ns
.PARAM t_b_485=4860.0ns
.PARAM t_b_486=4870.0215ns
.PARAM t_b_487=4880.0ns
.PARAM t_b_488=4890.022ns
.PARAM t_b_489=4900.0ns
.PARAM t_b_490=4910.0225ns
.PARAM t_b_491=4920.0ns
.PARAM t_b_492=4930.023ns
.PARAM t_b_493=4940.0ns
.PARAM t_b_494=4950.0235ns
.PARAM t_b_495=4960.0ns
.PARAM t_b_496=4970.024ns
.PARAM t_b_497=4980.0ns
.PARAM t_b_498=4990.0245ns
.PARAM t_b_499=5000.0ns
.PARAM t_b_500=5010.025ns
.PARAM t_b_501=5020.0ns
.PARAM t_b_502=5030.0255ns
.PARAM t_b_503=5040.0ns
.PARAM t_b_504=5050.026ns
.PARAM t_b_505=5060.0ns
.PARAM t_b_506=5070.0265ns
.PARAM t_b_507=5080.0ns
.PARAM t_b_508=5090.027ns
.PARAM t_b_509=5100.0ns
.PARAM t_b_510=5110.0275ns
.PARAM t_b_511=5120.0ns
.PARAM t_b_512=5130.028ns
.PARAM t_b_513=5140.0ns
.PARAM t_b_514=5150.0285ns
.PARAM t_b_515=5160.0ns
.PARAM t_b_516=5170.029ns
.PARAM t_b_517=5180.0ns
.PARAM t_b_518=5190.0295ns
.PARAM t_b_519=5200.0ns
.PARAM t_b_520=5210.03ns
.PARAM t_b_521=5220.0ns
.PARAM t_b_522=5230.0305ns
.PARAM t_b_523=5240.0ns
.PARAM t_b_524=5250.031ns
.PARAM t_b_525=5260.0ns
.PARAM t_b_526=5270.0315ns
.PARAM t_b_527=5280.0ns
.PARAM t_b_528=5290.032ns
.PARAM t_b_529=5300.0ns
.PARAM t_b_530=5310.0325ns
.PARAM t_b_531=5320.0ns
.PARAM t_b_532=5330.033ns
.PARAM t_b_533=5340.0ns
.PARAM t_b_534=5350.0335ns
.PARAM t_b_535=5360.0ns
.PARAM t_b_536=5370.034ns
.PARAM t_b_537=5380.0ns
.PARAM t_b_538=5390.0345ns
.PARAM t_b_539=5400.0ns
.PARAM t_b_540=5410.035ns
.PARAM t_b_541=5420.0ns
.PARAM t_b_542=5430.0355ns
.PARAM t_b_543=5440.0ns
.PARAM t_b_544=5450.036ns
.PARAM t_b_545=5460.0ns
.PARAM t_b_546=5470.0365ns
.PARAM t_b_547=5480.0ns
.PARAM t_b_548=5490.037ns
.PARAM t_b_549=5500.0ns
.PARAM t_b_550=5510.0375ns
.PARAM t_b_551=5520.0ns
.PARAM t_b_552=5530.038ns
.PARAM t_b_553=5540.0ns
.PARAM t_b_554=5550.0385ns
.PARAM t_b_555=5560.0ns
.PARAM t_b_556=5570.039ns
.PARAM t_b_557=5580.0ns
.PARAM t_b_558=5590.0395ns
.PARAM t_b_559=5600.0ns
.PARAM t_b_560=5610.04ns
.PARAM t_b_561=5620.0ns
.PARAM t_b_562=5630.0405ns
.PARAM t_b_563=5640.0ns
.PARAM t_b_564=5650.041ns
.PARAM t_b_565=5660.0ns
.PARAM t_b_566=5670.0415ns
.PARAM t_b_567=5680.0ns
.PARAM t_b_568=5690.042ns
.PARAM t_b_569=5700.0ns
.PARAM t_b_570=5710.0425ns
.PARAM t_b_571=5720.0ns
.PARAM t_b_572=5730.043ns
.PARAM t_b_573=5740.0ns
.PARAM t_b_574=5750.0435ns
.PARAM t_b_575=5760.0ns
.PARAM t_b_576=5770.044ns
.PARAM t_b_577=5780.0ns
.PARAM t_b_578=5790.0445ns
.PARAM t_b_579=5800.0ns
.PARAM t_b_580=5810.045ns
.PARAM t_b_581=5820.0ns
.PARAM t_b_582=5830.0455ns
.PARAM t_b_583=5840.0ns
.PARAM t_b_584=5850.046ns
.PARAM t_b_585=5860.0ns
.PARAM t_b_586=5870.0465ns
.PARAM t_b_587=5880.0ns
.PARAM t_b_588=5890.047ns
.PARAM t_b_589=5900.0ns
.PARAM t_b_590=5910.0475ns
.PARAM t_b_591=5920.0ns
.PARAM t_b_592=5930.048ns
.PARAM t_b_593=5940.0ns
.PARAM t_b_594=5950.0485ns
.PARAM t_b_595=5960.0ns
.PARAM t_b_596=5970.049ns
.PARAM t_b_597=5980.0ns
.PARAM t_b_598=5990.0495ns
.PARAM t_b_599=6000.0ns
.PARAM t_b_600=6010.05ns
.PARAM t_b_601=6020.0ns
.PARAM t_b_602=6030.0505ns
.PARAM t_b_603=6040.0ns
.PARAM t_b_604=6050.051ns
.PARAM t_b_605=6060.0ns
.PARAM t_b_606=6070.0515ns
.PARAM t_b_607=6080.0ns
.PARAM t_b_608=6090.052ns
.PARAM t_b_609=6100.0ns
.PARAM t_b_610=6110.0525ns
.PARAM t_b_611=6120.0ns
.PARAM t_b_612=6130.053ns
.PARAM t_b_613=6140.0ns
.PARAM t_b_614=6150.0535ns
.PARAM t_b_615=6160.0ns
.PARAM t_b_616=6170.054ns
.PARAM t_b_617=6180.0ns
.PARAM t_b_618=6190.0545ns
.PARAM t_b_619=6200.0ns
.PARAM t_b_620=6210.055ns
.PARAM t_b_621=6220.0ns
.PARAM t_b_622=6230.0555ns
.PARAM t_b_623=6240.0ns
.PARAM t_b_624=6250.056ns
.PARAM t_b_625=6260.0ns
.PARAM t_b_626=6270.0565ns
.PARAM t_b_627=6280.0ns
.PARAM t_b_628=6290.057ns
.PARAM t_b_629=6300.0ns
.PARAM t_b_630=6310.0575ns
.PARAM t_b_631=6320.0ns
.PARAM t_b_632=6330.058ns
.PARAM t_b_633=6340.0ns
.PARAM t_b_634=6350.0585ns
.PARAM t_b_635=6360.0ns
.PARAM t_b_636=6370.059ns
.PARAM t_b_637=6380.0ns
.PARAM t_b_638=6390.0595ns
.PARAM t_b_639=6400.0ns
.PARAM t_b_640=6410.06ns
.PARAM t_b_641=6420.0ns
.PARAM t_b_642=6430.0605ns
.PARAM t_b_643=6440.0ns
.PARAM t_b_644=6450.061ns
.PARAM t_b_645=6460.0ns
.PARAM t_b_646=6470.0615ns
.PARAM t_b_647=6480.0ns
.PARAM t_b_648=6490.062ns
.PARAM t_b_649=6500.0ns
.PARAM t_b_650=6510.0625ns
.PARAM t_b_651=6520.0ns
.PARAM t_b_652=6530.063ns
.PARAM t_b_653=6540.0ns
.PARAM t_b_654=6550.0635ns
.PARAM t_b_655=6560.0ns
.PARAM t_b_656=6570.064ns
.PARAM t_b_657=6580.0ns
.PARAM t_b_658=6590.0645ns
.PARAM t_b_659=6600.0ns
.PARAM t_b_660=6610.065ns
.PARAM t_b_661=6620.0ns
.PARAM t_b_662=6630.0655ns
.PARAM t_b_663=6640.0ns
.PARAM t_b_664=6650.066ns
.PARAM t_b_665=6660.0ns
.PARAM t_b_666=6670.0665ns
.PARAM t_b_667=6680.0ns
.PARAM t_b_668=6690.067ns
.PARAM t_b_669=6700.0ns
.PARAM t_b_670=6710.0675ns
.PARAM t_b_671=6720.0ns
.PARAM t_b_672=6730.068ns
.PARAM t_b_673=6740.0ns
.PARAM t_b_674=6750.0685ns
.PARAM t_b_675=6760.0ns
.PARAM t_b_676=6770.069ns
.PARAM t_b_677=6780.0ns
.PARAM t_b_678=6790.0695ns
.PARAM t_b_679=6800.0ns
.PARAM t_b_680=6810.07ns
.PARAM t_b_681=6820.0ns
.PARAM t_b_682=6830.0705ns
.PARAM t_b_683=6840.0ns
.PARAM t_b_684=6850.071ns
.PARAM t_b_685=6860.0ns
.PARAM t_b_686=6870.0715ns
.PARAM t_b_687=6880.0ns
.PARAM t_b_688=6890.072ns
.PARAM t_b_689=6900.0ns
.PARAM t_b_690=6910.0725ns
.PARAM t_b_691=6920.0ns
.PARAM t_b_692=6930.073ns
.PARAM t_b_693=6940.0ns
.PARAM t_b_694=6950.0735ns
.PARAM t_b_695=6960.0ns
.PARAM t_b_696=6970.074ns
.PARAM t_b_697=6980.0ns
.PARAM t_b_698=6990.0745ns
.PARAM t_b_699=7000.0ns
.PARAM t_b_700=7010.075ns
.PARAM t_b_701=7020.0ns
.PARAM t_b_702=7030.0755ns
.PARAM t_b_703=7040.0ns
.PARAM t_b_704=7050.076ns
.PARAM t_b_705=7060.0ns
.PARAM t_b_706=7070.0765ns
.PARAM t_b_707=7080.0ns
.PARAM t_b_708=7090.077ns
.PARAM t_b_709=7100.0ns
.PARAM t_b_710=7110.0775ns
.PARAM t_b_711=7120.0ns
.PARAM t_b_712=7130.078ns
.PARAM t_b_713=7140.0ns
.PARAM t_b_714=7150.0785ns
.PARAM t_b_715=7160.0ns
.PARAM t_b_716=7170.079ns
.PARAM t_b_717=7180.0ns
.PARAM t_b_718=7190.0795ns
.PARAM t_b_719=7200.0ns
.PARAM t_b_720=7210.08ns
.PARAM t_b_721=7220.0ns
.PARAM t_b_722=7230.0805ns
.PARAM t_b_723=7240.0ns
.PARAM t_b_724=7250.081ns
.PARAM t_b_725=7260.0ns
.PARAM t_b_726=7270.0815ns
.PARAM t_b_727=7280.0ns
.PARAM t_b_728=7290.082ns
.PARAM t_b_729=7300.0ns
.PARAM t_b_730=7310.0825ns
.PARAM t_b_731=7320.0ns
.PARAM t_b_732=7330.083ns
.PARAM t_b_733=7340.0ns
.PARAM t_b_734=7350.0835ns
.PARAM t_b_735=7360.0ns
.PARAM t_b_736=7370.084ns
.PARAM t_b_737=7380.0ns
.PARAM t_b_738=7390.0845ns
.PARAM t_b_739=7400.0ns
.PARAM t_b_740=7410.085ns
.PARAM t_b_741=7420.0ns
.PARAM t_b_742=7430.0855ns
.PARAM t_b_743=7440.0ns
.PARAM t_b_744=7450.086ns
.PARAM t_b_745=7460.0ns
.PARAM t_b_746=7470.0865ns
.PARAM t_b_747=7480.0ns
.PARAM t_b_748=7490.087ns
.PARAM t_b_749=7500.0ns
.PARAM t_b_750=7510.0875ns
.PARAM t_b_751=7520.0ns
.PARAM t_b_752=7530.088ns
.PARAM t_b_753=7540.0ns
.PARAM t_b_754=7550.0885ns
.PARAM t_b_755=7560.0ns
.PARAM t_b_756=7570.089ns
.PARAM t_b_757=7580.0ns
.PARAM t_b_758=7590.0895ns
.PARAM t_b_759=7600.0ns
.PARAM t_b_760=7610.09ns
.PARAM t_b_761=7620.0ns
.PARAM t_b_762=7630.0905ns
.PARAM t_b_763=7640.0ns
.PARAM t_b_764=7650.091ns
.PARAM t_b_765=7660.0ns
.PARAM t_b_766=7670.0915ns
.PARAM t_b_767=7680.0ns
.PARAM t_b_768=7690.092ns
.PARAM t_b_769=7700.0ns
.PARAM t_b_770=7710.0925ns
.PARAM t_b_771=7720.0ns
.PARAM t_b_772=7730.093ns
.PARAM t_b_773=7740.0ns
.PARAM t_b_774=7750.0935ns
.PARAM t_b_775=7760.0ns
.PARAM t_b_776=7770.094ns
.PARAM t_b_777=7780.0ns
.PARAM t_b_778=7790.0945ns
.PARAM t_b_779=7800.0ns
.PARAM t_b_780=7810.095ns
.PARAM t_b_781=7820.0ns
.PARAM t_b_782=7830.0955ns
.PARAM t_b_783=7840.0ns
.PARAM t_b_784=7850.096ns
.PARAM t_b_785=7860.0ns
.PARAM t_b_786=7870.0965ns
.PARAM t_b_787=7880.0ns
.PARAM t_b_788=7890.097ns
.PARAM t_b_789=7900.0ns
.PARAM t_b_790=7910.0975ns
.PARAM t_b_791=7920.0ns
.PARAM t_b_792=7930.098ns
.PARAM t_b_793=7940.0ns
.PARAM t_b_794=7950.0985ns
.PARAM t_b_795=7960.0ns
.PARAM t_b_796=7970.099ns
.PARAM t_b_797=7980.0ns
.PARAM t_b_798=7990.0995ns
.PARAM t_b_799=8000.0ns



VINA Input_A GND PWL 0ns baseVal t_init0 baseVal 't_init0+slope' peakVal t_init1 peakVal 't_init1+slope' baseVal
+ t_a_0 peakVal 't_a_0+slope' baseVal
+ t_a_1 baseVal 't_a_1+slope' peakVal
+ t_a_2 peakVal 't_a_2+slope' baseVal
+ t_a_3 baseVal 't_a_3+slope' peakVal
+ t_a_4 peakVal 't_a_4+slope' baseVal
+ t_a_5 baseVal 't_a_5+slope' peakVal
+ t_a_6 peakVal 't_a_6+slope' baseVal
+ t_a_7 baseVal 't_a_7+slope' peakVal
+ t_a_8 peakVal 't_a_8+slope' baseVal
+ t_a_9 baseVal 't_a_9+slope' peakVal
+ t_a_10 peakVal 't_a_10+slope' baseVal
+ t_a_11 baseVal 't_a_11+slope' peakVal
+ t_a_12 peakVal 't_a_12+slope' baseVal
+ t_a_13 baseVal 't_a_13+slope' peakVal
+ t_a_14 peakVal 't_a_14+slope' baseVal
+ t_a_15 baseVal 't_a_15+slope' peakVal
+ t_a_16 peakVal 't_a_16+slope' baseVal
+ t_a_17 baseVal 't_a_17+slope' peakVal
+ t_a_18 peakVal 't_a_18+slope' baseVal
+ t_a_19 baseVal 't_a_19+slope' peakVal
+ t_a_20 peakVal 't_a_20+slope' baseVal
+ t_a_21 baseVal 't_a_21+slope' peakVal
+ t_a_22 peakVal 't_a_22+slope' baseVal
+ t_a_23 baseVal 't_a_23+slope' peakVal
+ t_a_24 peakVal 't_a_24+slope' baseVal
+ t_a_25 baseVal 't_a_25+slope' peakVal
+ t_a_26 peakVal 't_a_26+slope' baseVal
+ t_a_27 baseVal 't_a_27+slope' peakVal
+ t_a_28 peakVal 't_a_28+slope' baseVal
+ t_a_29 baseVal 't_a_29+slope' peakVal
+ t_a_30 peakVal 't_a_30+slope' baseVal
+ t_a_31 baseVal 't_a_31+slope' peakVal
+ t_a_32 peakVal 't_a_32+slope' baseVal
+ t_a_33 baseVal 't_a_33+slope' peakVal
+ t_a_34 peakVal 't_a_34+slope' baseVal
+ t_a_35 baseVal 't_a_35+slope' peakVal
+ t_a_36 peakVal 't_a_36+slope' baseVal
+ t_a_37 baseVal 't_a_37+slope' peakVal
+ t_a_38 peakVal 't_a_38+slope' baseVal
+ t_a_39 baseVal 't_a_39+slope' peakVal
+ t_a_40 peakVal 't_a_40+slope' baseVal
+ t_a_41 baseVal 't_a_41+slope' peakVal
+ t_a_42 peakVal 't_a_42+slope' baseVal
+ t_a_43 baseVal 't_a_43+slope' peakVal
+ t_a_44 peakVal 't_a_44+slope' baseVal
+ t_a_45 baseVal 't_a_45+slope' peakVal
+ t_a_46 peakVal 't_a_46+slope' baseVal
+ t_a_47 baseVal 't_a_47+slope' peakVal
+ t_a_48 peakVal 't_a_48+slope' baseVal
+ t_a_49 baseVal 't_a_49+slope' peakVal
+ t_a_50 peakVal 't_a_50+slope' baseVal
+ t_a_51 baseVal 't_a_51+slope' peakVal
+ t_a_52 peakVal 't_a_52+slope' baseVal
+ t_a_53 baseVal 't_a_53+slope' peakVal
+ t_a_54 peakVal 't_a_54+slope' baseVal
+ t_a_55 baseVal 't_a_55+slope' peakVal
+ t_a_56 peakVal 't_a_56+slope' baseVal
+ t_a_57 baseVal 't_a_57+slope' peakVal
+ t_a_58 peakVal 't_a_58+slope' baseVal
+ t_a_59 baseVal 't_a_59+slope' peakVal
+ t_a_60 peakVal 't_a_60+slope' baseVal
+ t_a_61 baseVal 't_a_61+slope' peakVal
+ t_a_62 peakVal 't_a_62+slope' baseVal
+ t_a_63 baseVal 't_a_63+slope' peakVal
+ t_a_64 peakVal 't_a_64+slope' baseVal
+ t_a_65 baseVal 't_a_65+slope' peakVal
+ t_a_66 peakVal 't_a_66+slope' baseVal
+ t_a_67 baseVal 't_a_67+slope' peakVal
+ t_a_68 peakVal 't_a_68+slope' baseVal
+ t_a_69 baseVal 't_a_69+slope' peakVal
+ t_a_70 peakVal 't_a_70+slope' baseVal
+ t_a_71 baseVal 't_a_71+slope' peakVal
+ t_a_72 peakVal 't_a_72+slope' baseVal
+ t_a_73 baseVal 't_a_73+slope' peakVal
+ t_a_74 peakVal 't_a_74+slope' baseVal
+ t_a_75 baseVal 't_a_75+slope' peakVal
+ t_a_76 peakVal 't_a_76+slope' baseVal
+ t_a_77 baseVal 't_a_77+slope' peakVal
+ t_a_78 peakVal 't_a_78+slope' baseVal
+ t_a_79 baseVal 't_a_79+slope' peakVal
+ t_a_80 peakVal 't_a_80+slope' baseVal
+ t_a_81 baseVal 't_a_81+slope' peakVal
+ t_a_82 peakVal 't_a_82+slope' baseVal
+ t_a_83 baseVal 't_a_83+slope' peakVal
+ t_a_84 peakVal 't_a_84+slope' baseVal
+ t_a_85 baseVal 't_a_85+slope' peakVal
+ t_a_86 peakVal 't_a_86+slope' baseVal
+ t_a_87 baseVal 't_a_87+slope' peakVal
+ t_a_88 peakVal 't_a_88+slope' baseVal
+ t_a_89 baseVal 't_a_89+slope' peakVal
+ t_a_90 peakVal 't_a_90+slope' baseVal
+ t_a_91 baseVal 't_a_91+slope' peakVal
+ t_a_92 peakVal 't_a_92+slope' baseVal
+ t_a_93 baseVal 't_a_93+slope' peakVal
+ t_a_94 peakVal 't_a_94+slope' baseVal
+ t_a_95 baseVal 't_a_95+slope' peakVal
+ t_a_96 peakVal 't_a_96+slope' baseVal
+ t_a_97 baseVal 't_a_97+slope' peakVal
+ t_a_98 peakVal 't_a_98+slope' baseVal
+ t_a_99 baseVal 't_a_99+slope' peakVal
+ t_a_100 peakVal 't_a_100+slope' baseVal
+ t_a_101 baseVal 't_a_101+slope' peakVal
+ t_a_102 peakVal 't_a_102+slope' baseVal
+ t_a_103 baseVal 't_a_103+slope' peakVal
+ t_a_104 peakVal 't_a_104+slope' baseVal
+ t_a_105 baseVal 't_a_105+slope' peakVal
+ t_a_106 peakVal 't_a_106+slope' baseVal
+ t_a_107 baseVal 't_a_107+slope' peakVal
+ t_a_108 peakVal 't_a_108+slope' baseVal
+ t_a_109 baseVal 't_a_109+slope' peakVal
+ t_a_110 peakVal 't_a_110+slope' baseVal
+ t_a_111 baseVal 't_a_111+slope' peakVal
+ t_a_112 peakVal 't_a_112+slope' baseVal
+ t_a_113 baseVal 't_a_113+slope' peakVal
+ t_a_114 peakVal 't_a_114+slope' baseVal
+ t_a_115 baseVal 't_a_115+slope' peakVal
+ t_a_116 peakVal 't_a_116+slope' baseVal
+ t_a_117 baseVal 't_a_117+slope' peakVal
+ t_a_118 peakVal 't_a_118+slope' baseVal
+ t_a_119 baseVal 't_a_119+slope' peakVal
+ t_a_120 peakVal 't_a_120+slope' baseVal
+ t_a_121 baseVal 't_a_121+slope' peakVal
+ t_a_122 peakVal 't_a_122+slope' baseVal
+ t_a_123 baseVal 't_a_123+slope' peakVal
+ t_a_124 peakVal 't_a_124+slope' baseVal
+ t_a_125 baseVal 't_a_125+slope' peakVal
+ t_a_126 peakVal 't_a_126+slope' baseVal
+ t_a_127 baseVal 't_a_127+slope' peakVal
+ t_a_128 peakVal 't_a_128+slope' baseVal
+ t_a_129 baseVal 't_a_129+slope' peakVal
+ t_a_130 peakVal 't_a_130+slope' baseVal
+ t_a_131 baseVal 't_a_131+slope' peakVal
+ t_a_132 peakVal 't_a_132+slope' baseVal
+ t_a_133 baseVal 't_a_133+slope' peakVal
+ t_a_134 peakVal 't_a_134+slope' baseVal
+ t_a_135 baseVal 't_a_135+slope' peakVal
+ t_a_136 peakVal 't_a_136+slope' baseVal
+ t_a_137 baseVal 't_a_137+slope' peakVal
+ t_a_138 peakVal 't_a_138+slope' baseVal
+ t_a_139 baseVal 't_a_139+slope' peakVal
+ t_a_140 peakVal 't_a_140+slope' baseVal
+ t_a_141 baseVal 't_a_141+slope' peakVal
+ t_a_142 peakVal 't_a_142+slope' baseVal
+ t_a_143 baseVal 't_a_143+slope' peakVal
+ t_a_144 peakVal 't_a_144+slope' baseVal
+ t_a_145 baseVal 't_a_145+slope' peakVal
+ t_a_146 peakVal 't_a_146+slope' baseVal
+ t_a_147 baseVal 't_a_147+slope' peakVal
+ t_a_148 peakVal 't_a_148+slope' baseVal
+ t_a_149 baseVal 't_a_149+slope' peakVal
+ t_a_150 peakVal 't_a_150+slope' baseVal
+ t_a_151 baseVal 't_a_151+slope' peakVal
+ t_a_152 peakVal 't_a_152+slope' baseVal
+ t_a_153 baseVal 't_a_153+slope' peakVal
+ t_a_154 peakVal 't_a_154+slope' baseVal
+ t_a_155 baseVal 't_a_155+slope' peakVal
+ t_a_156 peakVal 't_a_156+slope' baseVal
+ t_a_157 baseVal 't_a_157+slope' peakVal
+ t_a_158 peakVal 't_a_158+slope' baseVal
+ t_a_159 baseVal 't_a_159+slope' peakVal
+ t_a_160 peakVal 't_a_160+slope' baseVal
+ t_a_161 baseVal 't_a_161+slope' peakVal
+ t_a_162 peakVal 't_a_162+slope' baseVal
+ t_a_163 baseVal 't_a_163+slope' peakVal
+ t_a_164 peakVal 't_a_164+slope' baseVal
+ t_a_165 baseVal 't_a_165+slope' peakVal
+ t_a_166 peakVal 't_a_166+slope' baseVal
+ t_a_167 baseVal 't_a_167+slope' peakVal
+ t_a_168 peakVal 't_a_168+slope' baseVal
+ t_a_169 baseVal 't_a_169+slope' peakVal
+ t_a_170 peakVal 't_a_170+slope' baseVal
+ t_a_171 baseVal 't_a_171+slope' peakVal
+ t_a_172 peakVal 't_a_172+slope' baseVal
+ t_a_173 baseVal 't_a_173+slope' peakVal
+ t_a_174 peakVal 't_a_174+slope' baseVal
+ t_a_175 baseVal 't_a_175+slope' peakVal
+ t_a_176 peakVal 't_a_176+slope' baseVal
+ t_a_177 baseVal 't_a_177+slope' peakVal
+ t_a_178 peakVal 't_a_178+slope' baseVal
+ t_a_179 baseVal 't_a_179+slope' peakVal
+ t_a_180 peakVal 't_a_180+slope' baseVal
+ t_a_181 baseVal 't_a_181+slope' peakVal
+ t_a_182 peakVal 't_a_182+slope' baseVal
+ t_a_183 baseVal 't_a_183+slope' peakVal
+ t_a_184 peakVal 't_a_184+slope' baseVal
+ t_a_185 baseVal 't_a_185+slope' peakVal
+ t_a_186 peakVal 't_a_186+slope' baseVal
+ t_a_187 baseVal 't_a_187+slope' peakVal
+ t_a_188 peakVal 't_a_188+slope' baseVal
+ t_a_189 baseVal 't_a_189+slope' peakVal
+ t_a_190 peakVal 't_a_190+slope' baseVal
+ t_a_191 baseVal 't_a_191+slope' peakVal
+ t_a_192 peakVal 't_a_192+slope' baseVal
+ t_a_193 baseVal 't_a_193+slope' peakVal
+ t_a_194 peakVal 't_a_194+slope' baseVal
+ t_a_195 baseVal 't_a_195+slope' peakVal
+ t_a_196 peakVal 't_a_196+slope' baseVal
+ t_a_197 baseVal 't_a_197+slope' peakVal
+ t_a_198 peakVal 't_a_198+slope' baseVal
+ t_a_199 baseVal 't_a_199+slope' peakVal
+ t_a_200 peakVal 't_a_200+slope' baseVal
+ t_a_201 baseVal 't_a_201+slope' peakVal
+ t_a_202 peakVal 't_a_202+slope' baseVal
+ t_a_203 baseVal 't_a_203+slope' peakVal
+ t_a_204 peakVal 't_a_204+slope' baseVal
+ t_a_205 baseVal 't_a_205+slope' peakVal
+ t_a_206 peakVal 't_a_206+slope' baseVal
+ t_a_207 baseVal 't_a_207+slope' peakVal
+ t_a_208 peakVal 't_a_208+slope' baseVal
+ t_a_209 baseVal 't_a_209+slope' peakVal
+ t_a_210 peakVal 't_a_210+slope' baseVal
+ t_a_211 baseVal 't_a_211+slope' peakVal
+ t_a_212 peakVal 't_a_212+slope' baseVal
+ t_a_213 baseVal 't_a_213+slope' peakVal
+ t_a_214 peakVal 't_a_214+slope' baseVal
+ t_a_215 baseVal 't_a_215+slope' peakVal
+ t_a_216 peakVal 't_a_216+slope' baseVal
+ t_a_217 baseVal 't_a_217+slope' peakVal
+ t_a_218 peakVal 't_a_218+slope' baseVal
+ t_a_219 baseVal 't_a_219+slope' peakVal
+ t_a_220 peakVal 't_a_220+slope' baseVal
+ t_a_221 baseVal 't_a_221+slope' peakVal
+ t_a_222 peakVal 't_a_222+slope' baseVal
+ t_a_223 baseVal 't_a_223+slope' peakVal
+ t_a_224 peakVal 't_a_224+slope' baseVal
+ t_a_225 baseVal 't_a_225+slope' peakVal
+ t_a_226 peakVal 't_a_226+slope' baseVal
+ t_a_227 baseVal 't_a_227+slope' peakVal
+ t_a_228 peakVal 't_a_228+slope' baseVal
+ t_a_229 baseVal 't_a_229+slope' peakVal
+ t_a_230 peakVal 't_a_230+slope' baseVal
+ t_a_231 baseVal 't_a_231+slope' peakVal
+ t_a_232 peakVal 't_a_232+slope' baseVal
+ t_a_233 baseVal 't_a_233+slope' peakVal
+ t_a_234 peakVal 't_a_234+slope' baseVal
+ t_a_235 baseVal 't_a_235+slope' peakVal
+ t_a_236 peakVal 't_a_236+slope' baseVal
+ t_a_237 baseVal 't_a_237+slope' peakVal
+ t_a_238 peakVal 't_a_238+slope' baseVal
+ t_a_239 baseVal 't_a_239+slope' peakVal
+ t_a_240 peakVal 't_a_240+slope' baseVal
+ t_a_241 baseVal 't_a_241+slope' peakVal
+ t_a_242 peakVal 't_a_242+slope' baseVal
+ t_a_243 baseVal 't_a_243+slope' peakVal
+ t_a_244 peakVal 't_a_244+slope' baseVal
+ t_a_245 baseVal 't_a_245+slope' peakVal
+ t_a_246 peakVal 't_a_246+slope' baseVal
+ t_a_247 baseVal 't_a_247+slope' peakVal
+ t_a_248 peakVal 't_a_248+slope' baseVal
+ t_a_249 baseVal 't_a_249+slope' peakVal
+ t_a_250 peakVal 't_a_250+slope' baseVal
+ t_a_251 baseVal 't_a_251+slope' peakVal
+ t_a_252 peakVal 't_a_252+slope' baseVal
+ t_a_253 baseVal 't_a_253+slope' peakVal
+ t_a_254 peakVal 't_a_254+slope' baseVal
+ t_a_255 baseVal 't_a_255+slope' peakVal
+ t_a_256 peakVal 't_a_256+slope' baseVal
+ t_a_257 baseVal 't_a_257+slope' peakVal
+ t_a_258 peakVal 't_a_258+slope' baseVal
+ t_a_259 baseVal 't_a_259+slope' peakVal
+ t_a_260 peakVal 't_a_260+slope' baseVal
+ t_a_261 baseVal 't_a_261+slope' peakVal
+ t_a_262 peakVal 't_a_262+slope' baseVal
+ t_a_263 baseVal 't_a_263+slope' peakVal
+ t_a_264 peakVal 't_a_264+slope' baseVal
+ t_a_265 baseVal 't_a_265+slope' peakVal
+ t_a_266 peakVal 't_a_266+slope' baseVal
+ t_a_267 baseVal 't_a_267+slope' peakVal
+ t_a_268 peakVal 't_a_268+slope' baseVal
+ t_a_269 baseVal 't_a_269+slope' peakVal
+ t_a_270 peakVal 't_a_270+slope' baseVal
+ t_a_271 baseVal 't_a_271+slope' peakVal
+ t_a_272 peakVal 't_a_272+slope' baseVal
+ t_a_273 baseVal 't_a_273+slope' peakVal
+ t_a_274 peakVal 't_a_274+slope' baseVal
+ t_a_275 baseVal 't_a_275+slope' peakVal
+ t_a_276 peakVal 't_a_276+slope' baseVal
+ t_a_277 baseVal 't_a_277+slope' peakVal
+ t_a_278 peakVal 't_a_278+slope' baseVal
+ t_a_279 baseVal 't_a_279+slope' peakVal
+ t_a_280 peakVal 't_a_280+slope' baseVal
+ t_a_281 baseVal 't_a_281+slope' peakVal
+ t_a_282 peakVal 't_a_282+slope' baseVal
+ t_a_283 baseVal 't_a_283+slope' peakVal
+ t_a_284 peakVal 't_a_284+slope' baseVal
+ t_a_285 baseVal 't_a_285+slope' peakVal
+ t_a_286 peakVal 't_a_286+slope' baseVal
+ t_a_287 baseVal 't_a_287+slope' peakVal
+ t_a_288 peakVal 't_a_288+slope' baseVal
+ t_a_289 baseVal 't_a_289+slope' peakVal
+ t_a_290 peakVal 't_a_290+slope' baseVal
+ t_a_291 baseVal 't_a_291+slope' peakVal
+ t_a_292 peakVal 't_a_292+slope' baseVal
+ t_a_293 baseVal 't_a_293+slope' peakVal
+ t_a_294 peakVal 't_a_294+slope' baseVal
+ t_a_295 baseVal 't_a_295+slope' peakVal
+ t_a_296 peakVal 't_a_296+slope' baseVal
+ t_a_297 baseVal 't_a_297+slope' peakVal
+ t_a_298 peakVal 't_a_298+slope' baseVal
+ t_a_299 baseVal 't_a_299+slope' peakVal
+ t_a_300 peakVal 't_a_300+slope' baseVal
+ t_a_301 baseVal 't_a_301+slope' peakVal
+ t_a_302 peakVal 't_a_302+slope' baseVal
+ t_a_303 baseVal 't_a_303+slope' peakVal
+ t_a_304 peakVal 't_a_304+slope' baseVal
+ t_a_305 baseVal 't_a_305+slope' peakVal
+ t_a_306 peakVal 't_a_306+slope' baseVal
+ t_a_307 baseVal 't_a_307+slope' peakVal
+ t_a_308 peakVal 't_a_308+slope' baseVal
+ t_a_309 baseVal 't_a_309+slope' peakVal
+ t_a_310 peakVal 't_a_310+slope' baseVal
+ t_a_311 baseVal 't_a_311+slope' peakVal
+ t_a_312 peakVal 't_a_312+slope' baseVal
+ t_a_313 baseVal 't_a_313+slope' peakVal
+ t_a_314 peakVal 't_a_314+slope' baseVal
+ t_a_315 baseVal 't_a_315+slope' peakVal
+ t_a_316 peakVal 't_a_316+slope' baseVal
+ t_a_317 baseVal 't_a_317+slope' peakVal
+ t_a_318 peakVal 't_a_318+slope' baseVal
+ t_a_319 baseVal 't_a_319+slope' peakVal
+ t_a_320 peakVal 't_a_320+slope' baseVal
+ t_a_321 baseVal 't_a_321+slope' peakVal
+ t_a_322 peakVal 't_a_322+slope' baseVal
+ t_a_323 baseVal 't_a_323+slope' peakVal
+ t_a_324 peakVal 't_a_324+slope' baseVal
+ t_a_325 baseVal 't_a_325+slope' peakVal
+ t_a_326 peakVal 't_a_326+slope' baseVal
+ t_a_327 baseVal 't_a_327+slope' peakVal
+ t_a_328 peakVal 't_a_328+slope' baseVal
+ t_a_329 baseVal 't_a_329+slope' peakVal
+ t_a_330 peakVal 't_a_330+slope' baseVal
+ t_a_331 baseVal 't_a_331+slope' peakVal
+ t_a_332 peakVal 't_a_332+slope' baseVal
+ t_a_333 baseVal 't_a_333+slope' peakVal
+ t_a_334 peakVal 't_a_334+slope' baseVal
+ t_a_335 baseVal 't_a_335+slope' peakVal
+ t_a_336 peakVal 't_a_336+slope' baseVal
+ t_a_337 baseVal 't_a_337+slope' peakVal
+ t_a_338 peakVal 't_a_338+slope' baseVal
+ t_a_339 baseVal 't_a_339+slope' peakVal
+ t_a_340 peakVal 't_a_340+slope' baseVal
+ t_a_341 baseVal 't_a_341+slope' peakVal
+ t_a_342 peakVal 't_a_342+slope' baseVal
+ t_a_343 baseVal 't_a_343+slope' peakVal
+ t_a_344 peakVal 't_a_344+slope' baseVal
+ t_a_345 baseVal 't_a_345+slope' peakVal
+ t_a_346 peakVal 't_a_346+slope' baseVal
+ t_a_347 baseVal 't_a_347+slope' peakVal
+ t_a_348 peakVal 't_a_348+slope' baseVal
+ t_a_349 baseVal 't_a_349+slope' peakVal
+ t_a_350 peakVal 't_a_350+slope' baseVal
+ t_a_351 baseVal 't_a_351+slope' peakVal
+ t_a_352 peakVal 't_a_352+slope' baseVal
+ t_a_353 baseVal 't_a_353+slope' peakVal
+ t_a_354 peakVal 't_a_354+slope' baseVal
+ t_a_355 baseVal 't_a_355+slope' peakVal
+ t_a_356 peakVal 't_a_356+slope' baseVal
+ t_a_357 baseVal 't_a_357+slope' peakVal
+ t_a_358 peakVal 't_a_358+slope' baseVal
+ t_a_359 baseVal 't_a_359+slope' peakVal
+ t_a_360 peakVal 't_a_360+slope' baseVal
+ t_a_361 baseVal 't_a_361+slope' peakVal
+ t_a_362 peakVal 't_a_362+slope' baseVal
+ t_a_363 baseVal 't_a_363+slope' peakVal
+ t_a_364 peakVal 't_a_364+slope' baseVal
+ t_a_365 baseVal 't_a_365+slope' peakVal
+ t_a_366 peakVal 't_a_366+slope' baseVal
+ t_a_367 baseVal 't_a_367+slope' peakVal
+ t_a_368 peakVal 't_a_368+slope' baseVal
+ t_a_369 baseVal 't_a_369+slope' peakVal
+ t_a_370 peakVal 't_a_370+slope' baseVal
+ t_a_371 baseVal 't_a_371+slope' peakVal
+ t_a_372 peakVal 't_a_372+slope' baseVal
+ t_a_373 baseVal 't_a_373+slope' peakVal
+ t_a_374 peakVal 't_a_374+slope' baseVal
+ t_a_375 baseVal 't_a_375+slope' peakVal
+ t_a_376 peakVal 't_a_376+slope' baseVal
+ t_a_377 baseVal 't_a_377+slope' peakVal
+ t_a_378 peakVal 't_a_378+slope' baseVal
+ t_a_379 baseVal 't_a_379+slope' peakVal
+ t_a_380 peakVal 't_a_380+slope' baseVal
+ t_a_381 baseVal 't_a_381+slope' peakVal
+ t_a_382 peakVal 't_a_382+slope' baseVal
+ t_a_383 baseVal 't_a_383+slope' peakVal
+ t_a_384 peakVal 't_a_384+slope' baseVal
+ t_a_385 baseVal 't_a_385+slope' peakVal
+ t_a_386 peakVal 't_a_386+slope' baseVal
+ t_a_387 baseVal 't_a_387+slope' peakVal
+ t_a_388 peakVal 't_a_388+slope' baseVal
+ t_a_389 baseVal 't_a_389+slope' peakVal
+ t_a_390 peakVal 't_a_390+slope' baseVal
+ t_a_391 baseVal 't_a_391+slope' peakVal
+ t_a_392 peakVal 't_a_392+slope' baseVal
+ t_a_393 baseVal 't_a_393+slope' peakVal
+ t_a_394 peakVal 't_a_394+slope' baseVal
+ t_a_395 baseVal 't_a_395+slope' peakVal
+ t_a_396 peakVal 't_a_396+slope' baseVal
+ t_a_397 baseVal 't_a_397+slope' peakVal
+ t_a_398 peakVal 't_a_398+slope' baseVal
+ t_a_399 baseVal 't_a_399+slope' peakVal
+ t_a_400 peakVal 't_a_400+slope' baseVal
+ t_a_401 baseVal 't_a_401+slope' peakVal
+ t_a_402 peakVal 't_a_402+slope' baseVal
+ t_a_403 baseVal 't_a_403+slope' peakVal
+ t_a_404 peakVal 't_a_404+slope' baseVal
+ t_a_405 baseVal 't_a_405+slope' peakVal
+ t_a_406 peakVal 't_a_406+slope' baseVal
+ t_a_407 baseVal 't_a_407+slope' peakVal
+ t_a_408 peakVal 't_a_408+slope' baseVal
+ t_a_409 baseVal 't_a_409+slope' peakVal
+ t_a_410 peakVal 't_a_410+slope' baseVal
+ t_a_411 baseVal 't_a_411+slope' peakVal
+ t_a_412 peakVal 't_a_412+slope' baseVal
+ t_a_413 baseVal 't_a_413+slope' peakVal
+ t_a_414 peakVal 't_a_414+slope' baseVal
+ t_a_415 baseVal 't_a_415+slope' peakVal
+ t_a_416 peakVal 't_a_416+slope' baseVal
+ t_a_417 baseVal 't_a_417+slope' peakVal
+ t_a_418 peakVal 't_a_418+slope' baseVal
+ t_a_419 baseVal 't_a_419+slope' peakVal
+ t_a_420 peakVal 't_a_420+slope' baseVal
+ t_a_421 baseVal 't_a_421+slope' peakVal
+ t_a_422 peakVal 't_a_422+slope' baseVal
+ t_a_423 baseVal 't_a_423+slope' peakVal
+ t_a_424 peakVal 't_a_424+slope' baseVal
+ t_a_425 baseVal 't_a_425+slope' peakVal
+ t_a_426 peakVal 't_a_426+slope' baseVal
+ t_a_427 baseVal 't_a_427+slope' peakVal
+ t_a_428 peakVal 't_a_428+slope' baseVal
+ t_a_429 baseVal 't_a_429+slope' peakVal
+ t_a_430 peakVal 't_a_430+slope' baseVal
+ t_a_431 baseVal 't_a_431+slope' peakVal
+ t_a_432 peakVal 't_a_432+slope' baseVal
+ t_a_433 baseVal 't_a_433+slope' peakVal
+ t_a_434 peakVal 't_a_434+slope' baseVal
+ t_a_435 baseVal 't_a_435+slope' peakVal
+ t_a_436 peakVal 't_a_436+slope' baseVal
+ t_a_437 baseVal 't_a_437+slope' peakVal
+ t_a_438 peakVal 't_a_438+slope' baseVal
+ t_a_439 baseVal 't_a_439+slope' peakVal
+ t_a_440 peakVal 't_a_440+slope' baseVal
+ t_a_441 baseVal 't_a_441+slope' peakVal
+ t_a_442 peakVal 't_a_442+slope' baseVal
+ t_a_443 baseVal 't_a_443+slope' peakVal
+ t_a_444 peakVal 't_a_444+slope' baseVal
+ t_a_445 baseVal 't_a_445+slope' peakVal
+ t_a_446 peakVal 't_a_446+slope' baseVal
+ t_a_447 baseVal 't_a_447+slope' peakVal
+ t_a_448 peakVal 't_a_448+slope' baseVal
+ t_a_449 baseVal 't_a_449+slope' peakVal
+ t_a_450 peakVal 't_a_450+slope' baseVal
+ t_a_451 baseVal 't_a_451+slope' peakVal
+ t_a_452 peakVal 't_a_452+slope' baseVal
+ t_a_453 baseVal 't_a_453+slope' peakVal
+ t_a_454 peakVal 't_a_454+slope' baseVal
+ t_a_455 baseVal 't_a_455+slope' peakVal
+ t_a_456 peakVal 't_a_456+slope' baseVal
+ t_a_457 baseVal 't_a_457+slope' peakVal
+ t_a_458 peakVal 't_a_458+slope' baseVal
+ t_a_459 baseVal 't_a_459+slope' peakVal
+ t_a_460 peakVal 't_a_460+slope' baseVal
+ t_a_461 baseVal 't_a_461+slope' peakVal
+ t_a_462 peakVal 't_a_462+slope' baseVal
+ t_a_463 baseVal 't_a_463+slope' peakVal
+ t_a_464 peakVal 't_a_464+slope' baseVal
+ t_a_465 baseVal 't_a_465+slope' peakVal
+ t_a_466 peakVal 't_a_466+slope' baseVal
+ t_a_467 baseVal 't_a_467+slope' peakVal
+ t_a_468 peakVal 't_a_468+slope' baseVal
+ t_a_469 baseVal 't_a_469+slope' peakVal
+ t_a_470 peakVal 't_a_470+slope' baseVal
+ t_a_471 baseVal 't_a_471+slope' peakVal
+ t_a_472 peakVal 't_a_472+slope' baseVal
+ t_a_473 baseVal 't_a_473+slope' peakVal
+ t_a_474 peakVal 't_a_474+slope' baseVal
+ t_a_475 baseVal 't_a_475+slope' peakVal
+ t_a_476 peakVal 't_a_476+slope' baseVal
+ t_a_477 baseVal 't_a_477+slope' peakVal
+ t_a_478 peakVal 't_a_478+slope' baseVal
+ t_a_479 baseVal 't_a_479+slope' peakVal
+ t_a_480 peakVal 't_a_480+slope' baseVal
+ t_a_481 baseVal 't_a_481+slope' peakVal
+ t_a_482 peakVal 't_a_482+slope' baseVal
+ t_a_483 baseVal 't_a_483+slope' peakVal
+ t_a_484 peakVal 't_a_484+slope' baseVal
+ t_a_485 baseVal 't_a_485+slope' peakVal
+ t_a_486 peakVal 't_a_486+slope' baseVal
+ t_a_487 baseVal 't_a_487+slope' peakVal
+ t_a_488 peakVal 't_a_488+slope' baseVal
+ t_a_489 baseVal 't_a_489+slope' peakVal
+ t_a_490 peakVal 't_a_490+slope' baseVal
+ t_a_491 baseVal 't_a_491+slope' peakVal
+ t_a_492 peakVal 't_a_492+slope' baseVal
+ t_a_493 baseVal 't_a_493+slope' peakVal
+ t_a_494 peakVal 't_a_494+slope' baseVal
+ t_a_495 baseVal 't_a_495+slope' peakVal
+ t_a_496 peakVal 't_a_496+slope' baseVal
+ t_a_497 baseVal 't_a_497+slope' peakVal
+ t_a_498 peakVal 't_a_498+slope' baseVal
+ t_a_499 baseVal 't_a_499+slope' peakVal
+ t_a_500 peakVal 't_a_500+slope' baseVal
+ t_a_501 baseVal 't_a_501+slope' peakVal
+ t_a_502 peakVal 't_a_502+slope' baseVal
+ t_a_503 baseVal 't_a_503+slope' peakVal
+ t_a_504 peakVal 't_a_504+slope' baseVal
+ t_a_505 baseVal 't_a_505+slope' peakVal
+ t_a_506 peakVal 't_a_506+slope' baseVal
+ t_a_507 baseVal 't_a_507+slope' peakVal
+ t_a_508 peakVal 't_a_508+slope' baseVal
+ t_a_509 baseVal 't_a_509+slope' peakVal
+ t_a_510 peakVal 't_a_510+slope' baseVal
+ t_a_511 baseVal 't_a_511+slope' peakVal
+ t_a_512 peakVal 't_a_512+slope' baseVal
+ t_a_513 baseVal 't_a_513+slope' peakVal
+ t_a_514 peakVal 't_a_514+slope' baseVal
+ t_a_515 baseVal 't_a_515+slope' peakVal
+ t_a_516 peakVal 't_a_516+slope' baseVal
+ t_a_517 baseVal 't_a_517+slope' peakVal
+ t_a_518 peakVal 't_a_518+slope' baseVal
+ t_a_519 baseVal 't_a_519+slope' peakVal
+ t_a_520 peakVal 't_a_520+slope' baseVal
+ t_a_521 baseVal 't_a_521+slope' peakVal
+ t_a_522 peakVal 't_a_522+slope' baseVal
+ t_a_523 baseVal 't_a_523+slope' peakVal
+ t_a_524 peakVal 't_a_524+slope' baseVal
+ t_a_525 baseVal 't_a_525+slope' peakVal
+ t_a_526 peakVal 't_a_526+slope' baseVal
+ t_a_527 baseVal 't_a_527+slope' peakVal
+ t_a_528 peakVal 't_a_528+slope' baseVal
+ t_a_529 baseVal 't_a_529+slope' peakVal
+ t_a_530 peakVal 't_a_530+slope' baseVal
+ t_a_531 baseVal 't_a_531+slope' peakVal
+ t_a_532 peakVal 't_a_532+slope' baseVal
+ t_a_533 baseVal 't_a_533+slope' peakVal
+ t_a_534 peakVal 't_a_534+slope' baseVal
+ t_a_535 baseVal 't_a_535+slope' peakVal
+ t_a_536 peakVal 't_a_536+slope' baseVal
+ t_a_537 baseVal 't_a_537+slope' peakVal
+ t_a_538 peakVal 't_a_538+slope' baseVal
+ t_a_539 baseVal 't_a_539+slope' peakVal
+ t_a_540 peakVal 't_a_540+slope' baseVal
+ t_a_541 baseVal 't_a_541+slope' peakVal
+ t_a_542 peakVal 't_a_542+slope' baseVal
+ t_a_543 baseVal 't_a_543+slope' peakVal
+ t_a_544 peakVal 't_a_544+slope' baseVal
+ t_a_545 baseVal 't_a_545+slope' peakVal
+ t_a_546 peakVal 't_a_546+slope' baseVal
+ t_a_547 baseVal 't_a_547+slope' peakVal
+ t_a_548 peakVal 't_a_548+slope' baseVal
+ t_a_549 baseVal 't_a_549+slope' peakVal
+ t_a_550 peakVal 't_a_550+slope' baseVal
+ t_a_551 baseVal 't_a_551+slope' peakVal
+ t_a_552 peakVal 't_a_552+slope' baseVal
+ t_a_553 baseVal 't_a_553+slope' peakVal
+ t_a_554 peakVal 't_a_554+slope' baseVal
+ t_a_555 baseVal 't_a_555+slope' peakVal
+ t_a_556 peakVal 't_a_556+slope' baseVal
+ t_a_557 baseVal 't_a_557+slope' peakVal
+ t_a_558 peakVal 't_a_558+slope' baseVal
+ t_a_559 baseVal 't_a_559+slope' peakVal
+ t_a_560 peakVal 't_a_560+slope' baseVal
+ t_a_561 baseVal 't_a_561+slope' peakVal
+ t_a_562 peakVal 't_a_562+slope' baseVal
+ t_a_563 baseVal 't_a_563+slope' peakVal
+ t_a_564 peakVal 't_a_564+slope' baseVal
+ t_a_565 baseVal 't_a_565+slope' peakVal
+ t_a_566 peakVal 't_a_566+slope' baseVal
+ t_a_567 baseVal 't_a_567+slope' peakVal
+ t_a_568 peakVal 't_a_568+slope' baseVal
+ t_a_569 baseVal 't_a_569+slope' peakVal
+ t_a_570 peakVal 't_a_570+slope' baseVal
+ t_a_571 baseVal 't_a_571+slope' peakVal
+ t_a_572 peakVal 't_a_572+slope' baseVal
+ t_a_573 baseVal 't_a_573+slope' peakVal
+ t_a_574 peakVal 't_a_574+slope' baseVal
+ t_a_575 baseVal 't_a_575+slope' peakVal
+ t_a_576 peakVal 't_a_576+slope' baseVal
+ t_a_577 baseVal 't_a_577+slope' peakVal
+ t_a_578 peakVal 't_a_578+slope' baseVal
+ t_a_579 baseVal 't_a_579+slope' peakVal
+ t_a_580 peakVal 't_a_580+slope' baseVal
+ t_a_581 baseVal 't_a_581+slope' peakVal
+ t_a_582 peakVal 't_a_582+slope' baseVal
+ t_a_583 baseVal 't_a_583+slope' peakVal
+ t_a_584 peakVal 't_a_584+slope' baseVal
+ t_a_585 baseVal 't_a_585+slope' peakVal
+ t_a_586 peakVal 't_a_586+slope' baseVal
+ t_a_587 baseVal 't_a_587+slope' peakVal
+ t_a_588 peakVal 't_a_588+slope' baseVal
+ t_a_589 baseVal 't_a_589+slope' peakVal
+ t_a_590 peakVal 't_a_590+slope' baseVal
+ t_a_591 baseVal 't_a_591+slope' peakVal
+ t_a_592 peakVal 't_a_592+slope' baseVal
+ t_a_593 baseVal 't_a_593+slope' peakVal
+ t_a_594 peakVal 't_a_594+slope' baseVal
+ t_a_595 baseVal 't_a_595+slope' peakVal
+ t_a_596 peakVal 't_a_596+slope' baseVal
+ t_a_597 baseVal 't_a_597+slope' peakVal
+ t_a_598 peakVal 't_a_598+slope' baseVal
+ t_a_599 baseVal 't_a_599+slope' peakVal
+ t_a_600 peakVal 't_a_600+slope' baseVal
+ t_a_601 baseVal 't_a_601+slope' peakVal
+ t_a_602 peakVal 't_a_602+slope' baseVal
+ t_a_603 baseVal 't_a_603+slope' peakVal
+ t_a_604 peakVal 't_a_604+slope' baseVal
+ t_a_605 baseVal 't_a_605+slope' peakVal
+ t_a_606 peakVal 't_a_606+slope' baseVal
+ t_a_607 baseVal 't_a_607+slope' peakVal
+ t_a_608 peakVal 't_a_608+slope' baseVal
+ t_a_609 baseVal 't_a_609+slope' peakVal
+ t_a_610 peakVal 't_a_610+slope' baseVal
+ t_a_611 baseVal 't_a_611+slope' peakVal
+ t_a_612 peakVal 't_a_612+slope' baseVal
+ t_a_613 baseVal 't_a_613+slope' peakVal
+ t_a_614 peakVal 't_a_614+slope' baseVal
+ t_a_615 baseVal 't_a_615+slope' peakVal
+ t_a_616 peakVal 't_a_616+slope' baseVal
+ t_a_617 baseVal 't_a_617+slope' peakVal
+ t_a_618 peakVal 't_a_618+slope' baseVal
+ t_a_619 baseVal 't_a_619+slope' peakVal
+ t_a_620 peakVal 't_a_620+slope' baseVal
+ t_a_621 baseVal 't_a_621+slope' peakVal
+ t_a_622 peakVal 't_a_622+slope' baseVal
+ t_a_623 baseVal 't_a_623+slope' peakVal
+ t_a_624 peakVal 't_a_624+slope' baseVal
+ t_a_625 baseVal 't_a_625+slope' peakVal
+ t_a_626 peakVal 't_a_626+slope' baseVal
+ t_a_627 baseVal 't_a_627+slope' peakVal
+ t_a_628 peakVal 't_a_628+slope' baseVal
+ t_a_629 baseVal 't_a_629+slope' peakVal
+ t_a_630 peakVal 't_a_630+slope' baseVal
+ t_a_631 baseVal 't_a_631+slope' peakVal
+ t_a_632 peakVal 't_a_632+slope' baseVal
+ t_a_633 baseVal 't_a_633+slope' peakVal
+ t_a_634 peakVal 't_a_634+slope' baseVal
+ t_a_635 baseVal 't_a_635+slope' peakVal
+ t_a_636 peakVal 't_a_636+slope' baseVal
+ t_a_637 baseVal 't_a_637+slope' peakVal
+ t_a_638 peakVal 't_a_638+slope' baseVal
+ t_a_639 baseVal 't_a_639+slope' peakVal
+ t_a_640 peakVal 't_a_640+slope' baseVal
+ t_a_641 baseVal 't_a_641+slope' peakVal
+ t_a_642 peakVal 't_a_642+slope' baseVal
+ t_a_643 baseVal 't_a_643+slope' peakVal
+ t_a_644 peakVal 't_a_644+slope' baseVal
+ t_a_645 baseVal 't_a_645+slope' peakVal
+ t_a_646 peakVal 't_a_646+slope' baseVal
+ t_a_647 baseVal 't_a_647+slope' peakVal
+ t_a_648 peakVal 't_a_648+slope' baseVal
+ t_a_649 baseVal 't_a_649+slope' peakVal
+ t_a_650 peakVal 't_a_650+slope' baseVal
+ t_a_651 baseVal 't_a_651+slope' peakVal
+ t_a_652 peakVal 't_a_652+slope' baseVal
+ t_a_653 baseVal 't_a_653+slope' peakVal
+ t_a_654 peakVal 't_a_654+slope' baseVal
+ t_a_655 baseVal 't_a_655+slope' peakVal
+ t_a_656 peakVal 't_a_656+slope' baseVal
+ t_a_657 baseVal 't_a_657+slope' peakVal
+ t_a_658 peakVal 't_a_658+slope' baseVal
+ t_a_659 baseVal 't_a_659+slope' peakVal
+ t_a_660 peakVal 't_a_660+slope' baseVal
+ t_a_661 baseVal 't_a_661+slope' peakVal
+ t_a_662 peakVal 't_a_662+slope' baseVal
+ t_a_663 baseVal 't_a_663+slope' peakVal
+ t_a_664 peakVal 't_a_664+slope' baseVal
+ t_a_665 baseVal 't_a_665+slope' peakVal
+ t_a_666 peakVal 't_a_666+slope' baseVal
+ t_a_667 baseVal 't_a_667+slope' peakVal
+ t_a_668 peakVal 't_a_668+slope' baseVal
+ t_a_669 baseVal 't_a_669+slope' peakVal
+ t_a_670 peakVal 't_a_670+slope' baseVal
+ t_a_671 baseVal 't_a_671+slope' peakVal
+ t_a_672 peakVal 't_a_672+slope' baseVal
+ t_a_673 baseVal 't_a_673+slope' peakVal
+ t_a_674 peakVal 't_a_674+slope' baseVal
+ t_a_675 baseVal 't_a_675+slope' peakVal
+ t_a_676 peakVal 't_a_676+slope' baseVal
+ t_a_677 baseVal 't_a_677+slope' peakVal
+ t_a_678 peakVal 't_a_678+slope' baseVal
+ t_a_679 baseVal 't_a_679+slope' peakVal
+ t_a_680 peakVal 't_a_680+slope' baseVal
+ t_a_681 baseVal 't_a_681+slope' peakVal
+ t_a_682 peakVal 't_a_682+slope' baseVal
+ t_a_683 baseVal 't_a_683+slope' peakVal
+ t_a_684 peakVal 't_a_684+slope' baseVal
+ t_a_685 baseVal 't_a_685+slope' peakVal
+ t_a_686 peakVal 't_a_686+slope' baseVal
+ t_a_687 baseVal 't_a_687+slope' peakVal
+ t_a_688 peakVal 't_a_688+slope' baseVal
+ t_a_689 baseVal 't_a_689+slope' peakVal
+ t_a_690 peakVal 't_a_690+slope' baseVal
+ t_a_691 baseVal 't_a_691+slope' peakVal
+ t_a_692 peakVal 't_a_692+slope' baseVal
+ t_a_693 baseVal 't_a_693+slope' peakVal
+ t_a_694 peakVal 't_a_694+slope' baseVal
+ t_a_695 baseVal 't_a_695+slope' peakVal
+ t_a_696 peakVal 't_a_696+slope' baseVal
+ t_a_697 baseVal 't_a_697+slope' peakVal
+ t_a_698 peakVal 't_a_698+slope' baseVal
+ t_a_699 baseVal 't_a_699+slope' peakVal
+ t_a_700 peakVal 't_a_700+slope' baseVal
+ t_a_701 baseVal 't_a_701+slope' peakVal
+ t_a_702 peakVal 't_a_702+slope' baseVal
+ t_a_703 baseVal 't_a_703+slope' peakVal
+ t_a_704 peakVal 't_a_704+slope' baseVal
+ t_a_705 baseVal 't_a_705+slope' peakVal
+ t_a_706 peakVal 't_a_706+slope' baseVal
+ t_a_707 baseVal 't_a_707+slope' peakVal
+ t_a_708 peakVal 't_a_708+slope' baseVal
+ t_a_709 baseVal 't_a_709+slope' peakVal
+ t_a_710 peakVal 't_a_710+slope' baseVal
+ t_a_711 baseVal 't_a_711+slope' peakVal
+ t_a_712 peakVal 't_a_712+slope' baseVal
+ t_a_713 baseVal 't_a_713+slope' peakVal
+ t_a_714 peakVal 't_a_714+slope' baseVal
+ t_a_715 baseVal 't_a_715+slope' peakVal
+ t_a_716 peakVal 't_a_716+slope' baseVal
+ t_a_717 baseVal 't_a_717+slope' peakVal
+ t_a_718 peakVal 't_a_718+slope' baseVal
+ t_a_719 baseVal 't_a_719+slope' peakVal
+ t_a_720 peakVal 't_a_720+slope' baseVal
+ t_a_721 baseVal 't_a_721+slope' peakVal
+ t_a_722 peakVal 't_a_722+slope' baseVal
+ t_a_723 baseVal 't_a_723+slope' peakVal
+ t_a_724 peakVal 't_a_724+slope' baseVal
+ t_a_725 baseVal 't_a_725+slope' peakVal
+ t_a_726 peakVal 't_a_726+slope' baseVal
+ t_a_727 baseVal 't_a_727+slope' peakVal
+ t_a_728 peakVal 't_a_728+slope' baseVal
+ t_a_729 baseVal 't_a_729+slope' peakVal
+ t_a_730 peakVal 't_a_730+slope' baseVal
+ t_a_731 baseVal 't_a_731+slope' peakVal
+ t_a_732 peakVal 't_a_732+slope' baseVal
+ t_a_733 baseVal 't_a_733+slope' peakVal
+ t_a_734 peakVal 't_a_734+slope' baseVal
+ t_a_735 baseVal 't_a_735+slope' peakVal
+ t_a_736 peakVal 't_a_736+slope' baseVal
+ t_a_737 baseVal 't_a_737+slope' peakVal
+ t_a_738 peakVal 't_a_738+slope' baseVal
+ t_a_739 baseVal 't_a_739+slope' peakVal
+ t_a_740 peakVal 't_a_740+slope' baseVal
+ t_a_741 baseVal 't_a_741+slope' peakVal
+ t_a_742 peakVal 't_a_742+slope' baseVal
+ t_a_743 baseVal 't_a_743+slope' peakVal
+ t_a_744 peakVal 't_a_744+slope' baseVal
+ t_a_745 baseVal 't_a_745+slope' peakVal
+ t_a_746 peakVal 't_a_746+slope' baseVal
+ t_a_747 baseVal 't_a_747+slope' peakVal
+ t_a_748 peakVal 't_a_748+slope' baseVal
+ t_a_749 baseVal 't_a_749+slope' peakVal
+ t_a_750 peakVal 't_a_750+slope' baseVal
+ t_a_751 baseVal 't_a_751+slope' peakVal
+ t_a_752 peakVal 't_a_752+slope' baseVal
+ t_a_753 baseVal 't_a_753+slope' peakVal
+ t_a_754 peakVal 't_a_754+slope' baseVal
+ t_a_755 baseVal 't_a_755+slope' peakVal
+ t_a_756 peakVal 't_a_756+slope' baseVal
+ t_a_757 baseVal 't_a_757+slope' peakVal
+ t_a_758 peakVal 't_a_758+slope' baseVal
+ t_a_759 baseVal 't_a_759+slope' peakVal
+ t_a_760 peakVal 't_a_760+slope' baseVal
+ t_a_761 baseVal 't_a_761+slope' peakVal
+ t_a_762 peakVal 't_a_762+slope' baseVal
+ t_a_763 baseVal 't_a_763+slope' peakVal
+ t_a_764 peakVal 't_a_764+slope' baseVal
+ t_a_765 baseVal 't_a_765+slope' peakVal
+ t_a_766 peakVal 't_a_766+slope' baseVal
+ t_a_767 baseVal 't_a_767+slope' peakVal
+ t_a_768 peakVal 't_a_768+slope' baseVal
+ t_a_769 baseVal 't_a_769+slope' peakVal
+ t_a_770 peakVal 't_a_770+slope' baseVal
+ t_a_771 baseVal 't_a_771+slope' peakVal
+ t_a_772 peakVal 't_a_772+slope' baseVal
+ t_a_773 baseVal 't_a_773+slope' peakVal
+ t_a_774 peakVal 't_a_774+slope' baseVal
+ t_a_775 baseVal 't_a_775+slope' peakVal
+ t_a_776 peakVal 't_a_776+slope' baseVal
+ t_a_777 baseVal 't_a_777+slope' peakVal
+ t_a_778 peakVal 't_a_778+slope' baseVal
+ t_a_779 baseVal 't_a_779+slope' peakVal
+ t_a_780 peakVal 't_a_780+slope' baseVal
+ t_a_781 baseVal 't_a_781+slope' peakVal
+ t_a_782 peakVal 't_a_782+slope' baseVal
+ t_a_783 baseVal 't_a_783+slope' peakVal
+ t_a_784 peakVal 't_a_784+slope' baseVal
+ t_a_785 baseVal 't_a_785+slope' peakVal
+ t_a_786 peakVal 't_a_786+slope' baseVal
+ t_a_787 baseVal 't_a_787+slope' peakVal
+ t_a_788 peakVal 't_a_788+slope' baseVal
+ t_a_789 baseVal 't_a_789+slope' peakVal
+ t_a_790 peakVal 't_a_790+slope' baseVal
+ t_a_791 baseVal 't_a_791+slope' peakVal
+ t_a_792 peakVal 't_a_792+slope' baseVal
+ t_a_793 baseVal 't_a_793+slope' peakVal
+ t_a_794 peakVal 't_a_794+slope' baseVal
+ t_a_795 baseVal 't_a_795+slope' peakVal
+ t_a_796 peakVal 't_a_796+slope' baseVal
+ t_a_797 baseVal 't_a_797+slope' peakVal
+ t_a_798 peakVal 't_a_798+slope' baseVal
+ t_a_799 baseVal 't_a_799+slope' peakVal



VINB Input_B GND PWL 0ns baseVal t_init0 baseVal 't_init0+slope' peakVal t_init1 peakVal 't_init1+slope' baseVal
+ t_b_0 peakVal 't_b_0+slope' baseVal
+ t_b_1 baseVal 't_b_1+slope' peakVal
+ t_b_2 peakVal 't_b_2+slope' baseVal
+ t_b_3 baseVal 't_b_3+slope' peakVal
+ t_b_4 peakVal 't_b_4+slope' baseVal
+ t_b_5 baseVal 't_b_5+slope' peakVal
+ t_b_6 peakVal 't_b_6+slope' baseVal
+ t_b_7 baseVal 't_b_7+slope' peakVal
+ t_b_8 peakVal 't_b_8+slope' baseVal
+ t_b_9 baseVal 't_b_9+slope' peakVal
+ t_b_10 peakVal 't_b_10+slope' baseVal
+ t_b_11 baseVal 't_b_11+slope' peakVal
+ t_b_12 peakVal 't_b_12+slope' baseVal
+ t_b_13 baseVal 't_b_13+slope' peakVal
+ t_b_14 peakVal 't_b_14+slope' baseVal
+ t_b_15 baseVal 't_b_15+slope' peakVal
+ t_b_16 peakVal 't_b_16+slope' baseVal
+ t_b_17 baseVal 't_b_17+slope' peakVal
+ t_b_18 peakVal 't_b_18+slope' baseVal
+ t_b_19 baseVal 't_b_19+slope' peakVal
+ t_b_20 peakVal 't_b_20+slope' baseVal
+ t_b_21 baseVal 't_b_21+slope' peakVal
+ t_b_22 peakVal 't_b_22+slope' baseVal
+ t_b_23 baseVal 't_b_23+slope' peakVal
+ t_b_24 peakVal 't_b_24+slope' baseVal
+ t_b_25 baseVal 't_b_25+slope' peakVal
+ t_b_26 peakVal 't_b_26+slope' baseVal
+ t_b_27 baseVal 't_b_27+slope' peakVal
+ t_b_28 peakVal 't_b_28+slope' baseVal
+ t_b_29 baseVal 't_b_29+slope' peakVal
+ t_b_30 peakVal 't_b_30+slope' baseVal
+ t_b_31 baseVal 't_b_31+slope' peakVal
+ t_b_32 peakVal 't_b_32+slope' baseVal
+ t_b_33 baseVal 't_b_33+slope' peakVal
+ t_b_34 peakVal 't_b_34+slope' baseVal
+ t_b_35 baseVal 't_b_35+slope' peakVal
+ t_b_36 peakVal 't_b_36+slope' baseVal
+ t_b_37 baseVal 't_b_37+slope' peakVal
+ t_b_38 peakVal 't_b_38+slope' baseVal
+ t_b_39 baseVal 't_b_39+slope' peakVal
+ t_b_40 peakVal 't_b_40+slope' baseVal
+ t_b_41 baseVal 't_b_41+slope' peakVal
+ t_b_42 peakVal 't_b_42+slope' baseVal
+ t_b_43 baseVal 't_b_43+slope' peakVal
+ t_b_44 peakVal 't_b_44+slope' baseVal
+ t_b_45 baseVal 't_b_45+slope' peakVal
+ t_b_46 peakVal 't_b_46+slope' baseVal
+ t_b_47 baseVal 't_b_47+slope' peakVal
+ t_b_48 peakVal 't_b_48+slope' baseVal
+ t_b_49 baseVal 't_b_49+slope' peakVal
+ t_b_50 peakVal 't_b_50+slope' baseVal
+ t_b_51 baseVal 't_b_51+slope' peakVal
+ t_b_52 peakVal 't_b_52+slope' baseVal
+ t_b_53 baseVal 't_b_53+slope' peakVal
+ t_b_54 peakVal 't_b_54+slope' baseVal
+ t_b_55 baseVal 't_b_55+slope' peakVal
+ t_b_56 peakVal 't_b_56+slope' baseVal
+ t_b_57 baseVal 't_b_57+slope' peakVal
+ t_b_58 peakVal 't_b_58+slope' baseVal
+ t_b_59 baseVal 't_b_59+slope' peakVal
+ t_b_60 peakVal 't_b_60+slope' baseVal
+ t_b_61 baseVal 't_b_61+slope' peakVal
+ t_b_62 peakVal 't_b_62+slope' baseVal
+ t_b_63 baseVal 't_b_63+slope' peakVal
+ t_b_64 peakVal 't_b_64+slope' baseVal
+ t_b_65 baseVal 't_b_65+slope' peakVal
+ t_b_66 peakVal 't_b_66+slope' baseVal
+ t_b_67 baseVal 't_b_67+slope' peakVal
+ t_b_68 peakVal 't_b_68+slope' baseVal
+ t_b_69 baseVal 't_b_69+slope' peakVal
+ t_b_70 peakVal 't_b_70+slope' baseVal
+ t_b_71 baseVal 't_b_71+slope' peakVal
+ t_b_72 peakVal 't_b_72+slope' baseVal
+ t_b_73 baseVal 't_b_73+slope' peakVal
+ t_b_74 peakVal 't_b_74+slope' baseVal
+ t_b_75 baseVal 't_b_75+slope' peakVal
+ t_b_76 peakVal 't_b_76+slope' baseVal
+ t_b_77 baseVal 't_b_77+slope' peakVal
+ t_b_78 peakVal 't_b_78+slope' baseVal
+ t_b_79 baseVal 't_b_79+slope' peakVal
+ t_b_80 peakVal 't_b_80+slope' baseVal
+ t_b_81 baseVal 't_b_81+slope' peakVal
+ t_b_82 peakVal 't_b_82+slope' baseVal
+ t_b_83 baseVal 't_b_83+slope' peakVal
+ t_b_84 peakVal 't_b_84+slope' baseVal
+ t_b_85 baseVal 't_b_85+slope' peakVal
+ t_b_86 peakVal 't_b_86+slope' baseVal
+ t_b_87 baseVal 't_b_87+slope' peakVal
+ t_b_88 peakVal 't_b_88+slope' baseVal
+ t_b_89 baseVal 't_b_89+slope' peakVal
+ t_b_90 peakVal 't_b_90+slope' baseVal
+ t_b_91 baseVal 't_b_91+slope' peakVal
+ t_b_92 peakVal 't_b_92+slope' baseVal
+ t_b_93 baseVal 't_b_93+slope' peakVal
+ t_b_94 peakVal 't_b_94+slope' baseVal
+ t_b_95 baseVal 't_b_95+slope' peakVal
+ t_b_96 peakVal 't_b_96+slope' baseVal
+ t_b_97 baseVal 't_b_97+slope' peakVal
+ t_b_98 peakVal 't_b_98+slope' baseVal
+ t_b_99 baseVal 't_b_99+slope' peakVal
+ t_b_100 peakVal 't_b_100+slope' baseVal
+ t_b_101 baseVal 't_b_101+slope' peakVal
+ t_b_102 peakVal 't_b_102+slope' baseVal
+ t_b_103 baseVal 't_b_103+slope' peakVal
+ t_b_104 peakVal 't_b_104+slope' baseVal
+ t_b_105 baseVal 't_b_105+slope' peakVal
+ t_b_106 peakVal 't_b_106+slope' baseVal
+ t_b_107 baseVal 't_b_107+slope' peakVal
+ t_b_108 peakVal 't_b_108+slope' baseVal
+ t_b_109 baseVal 't_b_109+slope' peakVal
+ t_b_110 peakVal 't_b_110+slope' baseVal
+ t_b_111 baseVal 't_b_111+slope' peakVal
+ t_b_112 peakVal 't_b_112+slope' baseVal
+ t_b_113 baseVal 't_b_113+slope' peakVal
+ t_b_114 peakVal 't_b_114+slope' baseVal
+ t_b_115 baseVal 't_b_115+slope' peakVal
+ t_b_116 peakVal 't_b_116+slope' baseVal
+ t_b_117 baseVal 't_b_117+slope' peakVal
+ t_b_118 peakVal 't_b_118+slope' baseVal
+ t_b_119 baseVal 't_b_119+slope' peakVal
+ t_b_120 peakVal 't_b_120+slope' baseVal
+ t_b_121 baseVal 't_b_121+slope' peakVal
+ t_b_122 peakVal 't_b_122+slope' baseVal
+ t_b_123 baseVal 't_b_123+slope' peakVal
+ t_b_124 peakVal 't_b_124+slope' baseVal
+ t_b_125 baseVal 't_b_125+slope' peakVal
+ t_b_126 peakVal 't_b_126+slope' baseVal
+ t_b_127 baseVal 't_b_127+slope' peakVal
+ t_b_128 peakVal 't_b_128+slope' baseVal
+ t_b_129 baseVal 't_b_129+slope' peakVal
+ t_b_130 peakVal 't_b_130+slope' baseVal
+ t_b_131 baseVal 't_b_131+slope' peakVal
+ t_b_132 peakVal 't_b_132+slope' baseVal
+ t_b_133 baseVal 't_b_133+slope' peakVal
+ t_b_134 peakVal 't_b_134+slope' baseVal
+ t_b_135 baseVal 't_b_135+slope' peakVal
+ t_b_136 peakVal 't_b_136+slope' baseVal
+ t_b_137 baseVal 't_b_137+slope' peakVal
+ t_b_138 peakVal 't_b_138+slope' baseVal
+ t_b_139 baseVal 't_b_139+slope' peakVal
+ t_b_140 peakVal 't_b_140+slope' baseVal
+ t_b_141 baseVal 't_b_141+slope' peakVal
+ t_b_142 peakVal 't_b_142+slope' baseVal
+ t_b_143 baseVal 't_b_143+slope' peakVal
+ t_b_144 peakVal 't_b_144+slope' baseVal
+ t_b_145 baseVal 't_b_145+slope' peakVal
+ t_b_146 peakVal 't_b_146+slope' baseVal
+ t_b_147 baseVal 't_b_147+slope' peakVal
+ t_b_148 peakVal 't_b_148+slope' baseVal
+ t_b_149 baseVal 't_b_149+slope' peakVal
+ t_b_150 peakVal 't_b_150+slope' baseVal
+ t_b_151 baseVal 't_b_151+slope' peakVal
+ t_b_152 peakVal 't_b_152+slope' baseVal
+ t_b_153 baseVal 't_b_153+slope' peakVal
+ t_b_154 peakVal 't_b_154+slope' baseVal
+ t_b_155 baseVal 't_b_155+slope' peakVal
+ t_b_156 peakVal 't_b_156+slope' baseVal
+ t_b_157 baseVal 't_b_157+slope' peakVal
+ t_b_158 peakVal 't_b_158+slope' baseVal
+ t_b_159 baseVal 't_b_159+slope' peakVal
+ t_b_160 peakVal 't_b_160+slope' baseVal
+ t_b_161 baseVal 't_b_161+slope' peakVal
+ t_b_162 peakVal 't_b_162+slope' baseVal
+ t_b_163 baseVal 't_b_163+slope' peakVal
+ t_b_164 peakVal 't_b_164+slope' baseVal
+ t_b_165 baseVal 't_b_165+slope' peakVal
+ t_b_166 peakVal 't_b_166+slope' baseVal
+ t_b_167 baseVal 't_b_167+slope' peakVal
+ t_b_168 peakVal 't_b_168+slope' baseVal
+ t_b_169 baseVal 't_b_169+slope' peakVal
+ t_b_170 peakVal 't_b_170+slope' baseVal
+ t_b_171 baseVal 't_b_171+slope' peakVal
+ t_b_172 peakVal 't_b_172+slope' baseVal
+ t_b_173 baseVal 't_b_173+slope' peakVal
+ t_b_174 peakVal 't_b_174+slope' baseVal
+ t_b_175 baseVal 't_b_175+slope' peakVal
+ t_b_176 peakVal 't_b_176+slope' baseVal
+ t_b_177 baseVal 't_b_177+slope' peakVal
+ t_b_178 peakVal 't_b_178+slope' baseVal
+ t_b_179 baseVal 't_b_179+slope' peakVal
+ t_b_180 peakVal 't_b_180+slope' baseVal
+ t_b_181 baseVal 't_b_181+slope' peakVal
+ t_b_182 peakVal 't_b_182+slope' baseVal
+ t_b_183 baseVal 't_b_183+slope' peakVal
+ t_b_184 peakVal 't_b_184+slope' baseVal
+ t_b_185 baseVal 't_b_185+slope' peakVal
+ t_b_186 peakVal 't_b_186+slope' baseVal
+ t_b_187 baseVal 't_b_187+slope' peakVal
+ t_b_188 peakVal 't_b_188+slope' baseVal
+ t_b_189 baseVal 't_b_189+slope' peakVal
+ t_b_190 peakVal 't_b_190+slope' baseVal
+ t_b_191 baseVal 't_b_191+slope' peakVal
+ t_b_192 peakVal 't_b_192+slope' baseVal
+ t_b_193 baseVal 't_b_193+slope' peakVal
+ t_b_194 peakVal 't_b_194+slope' baseVal
+ t_b_195 baseVal 't_b_195+slope' peakVal
+ t_b_196 peakVal 't_b_196+slope' baseVal
+ t_b_197 baseVal 't_b_197+slope' peakVal
+ t_b_198 peakVal 't_b_198+slope' baseVal
+ t_b_199 baseVal 't_b_199+slope' peakVal
+ t_b_200 peakVal 't_b_200+slope' baseVal
+ t_b_201 baseVal 't_b_201+slope' peakVal
+ t_b_202 peakVal 't_b_202+slope' baseVal
+ t_b_203 baseVal 't_b_203+slope' peakVal
+ t_b_204 peakVal 't_b_204+slope' baseVal
+ t_b_205 baseVal 't_b_205+slope' peakVal
+ t_b_206 peakVal 't_b_206+slope' baseVal
+ t_b_207 baseVal 't_b_207+slope' peakVal
+ t_b_208 peakVal 't_b_208+slope' baseVal
+ t_b_209 baseVal 't_b_209+slope' peakVal
+ t_b_210 peakVal 't_b_210+slope' baseVal
+ t_b_211 baseVal 't_b_211+slope' peakVal
+ t_b_212 peakVal 't_b_212+slope' baseVal
+ t_b_213 baseVal 't_b_213+slope' peakVal
+ t_b_214 peakVal 't_b_214+slope' baseVal
+ t_b_215 baseVal 't_b_215+slope' peakVal
+ t_b_216 peakVal 't_b_216+slope' baseVal
+ t_b_217 baseVal 't_b_217+slope' peakVal
+ t_b_218 peakVal 't_b_218+slope' baseVal
+ t_b_219 baseVal 't_b_219+slope' peakVal
+ t_b_220 peakVal 't_b_220+slope' baseVal
+ t_b_221 baseVal 't_b_221+slope' peakVal
+ t_b_222 peakVal 't_b_222+slope' baseVal
+ t_b_223 baseVal 't_b_223+slope' peakVal
+ t_b_224 peakVal 't_b_224+slope' baseVal
+ t_b_225 baseVal 't_b_225+slope' peakVal
+ t_b_226 peakVal 't_b_226+slope' baseVal
+ t_b_227 baseVal 't_b_227+slope' peakVal
+ t_b_228 peakVal 't_b_228+slope' baseVal
+ t_b_229 baseVal 't_b_229+slope' peakVal
+ t_b_230 peakVal 't_b_230+slope' baseVal
+ t_b_231 baseVal 't_b_231+slope' peakVal
+ t_b_232 peakVal 't_b_232+slope' baseVal
+ t_b_233 baseVal 't_b_233+slope' peakVal
+ t_b_234 peakVal 't_b_234+slope' baseVal
+ t_b_235 baseVal 't_b_235+slope' peakVal
+ t_b_236 peakVal 't_b_236+slope' baseVal
+ t_b_237 baseVal 't_b_237+slope' peakVal
+ t_b_238 peakVal 't_b_238+slope' baseVal
+ t_b_239 baseVal 't_b_239+slope' peakVal
+ t_b_240 peakVal 't_b_240+slope' baseVal
+ t_b_241 baseVal 't_b_241+slope' peakVal
+ t_b_242 peakVal 't_b_242+slope' baseVal
+ t_b_243 baseVal 't_b_243+slope' peakVal
+ t_b_244 peakVal 't_b_244+slope' baseVal
+ t_b_245 baseVal 't_b_245+slope' peakVal
+ t_b_246 peakVal 't_b_246+slope' baseVal
+ t_b_247 baseVal 't_b_247+slope' peakVal
+ t_b_248 peakVal 't_b_248+slope' baseVal
+ t_b_249 baseVal 't_b_249+slope' peakVal
+ t_b_250 peakVal 't_b_250+slope' baseVal
+ t_b_251 baseVal 't_b_251+slope' peakVal
+ t_b_252 peakVal 't_b_252+slope' baseVal
+ t_b_253 baseVal 't_b_253+slope' peakVal
+ t_b_254 peakVal 't_b_254+slope' baseVal
+ t_b_255 baseVal 't_b_255+slope' peakVal
+ t_b_256 peakVal 't_b_256+slope' baseVal
+ t_b_257 baseVal 't_b_257+slope' peakVal
+ t_b_258 peakVal 't_b_258+slope' baseVal
+ t_b_259 baseVal 't_b_259+slope' peakVal
+ t_b_260 peakVal 't_b_260+slope' baseVal
+ t_b_261 baseVal 't_b_261+slope' peakVal
+ t_b_262 peakVal 't_b_262+slope' baseVal
+ t_b_263 baseVal 't_b_263+slope' peakVal
+ t_b_264 peakVal 't_b_264+slope' baseVal
+ t_b_265 baseVal 't_b_265+slope' peakVal
+ t_b_266 peakVal 't_b_266+slope' baseVal
+ t_b_267 baseVal 't_b_267+slope' peakVal
+ t_b_268 peakVal 't_b_268+slope' baseVal
+ t_b_269 baseVal 't_b_269+slope' peakVal
+ t_b_270 peakVal 't_b_270+slope' baseVal
+ t_b_271 baseVal 't_b_271+slope' peakVal
+ t_b_272 peakVal 't_b_272+slope' baseVal
+ t_b_273 baseVal 't_b_273+slope' peakVal
+ t_b_274 peakVal 't_b_274+slope' baseVal
+ t_b_275 baseVal 't_b_275+slope' peakVal
+ t_b_276 peakVal 't_b_276+slope' baseVal
+ t_b_277 baseVal 't_b_277+slope' peakVal
+ t_b_278 peakVal 't_b_278+slope' baseVal
+ t_b_279 baseVal 't_b_279+slope' peakVal
+ t_b_280 peakVal 't_b_280+slope' baseVal
+ t_b_281 baseVal 't_b_281+slope' peakVal
+ t_b_282 peakVal 't_b_282+slope' baseVal
+ t_b_283 baseVal 't_b_283+slope' peakVal
+ t_b_284 peakVal 't_b_284+slope' baseVal
+ t_b_285 baseVal 't_b_285+slope' peakVal
+ t_b_286 peakVal 't_b_286+slope' baseVal
+ t_b_287 baseVal 't_b_287+slope' peakVal
+ t_b_288 peakVal 't_b_288+slope' baseVal
+ t_b_289 baseVal 't_b_289+slope' peakVal
+ t_b_290 peakVal 't_b_290+slope' baseVal
+ t_b_291 baseVal 't_b_291+slope' peakVal
+ t_b_292 peakVal 't_b_292+slope' baseVal
+ t_b_293 baseVal 't_b_293+slope' peakVal
+ t_b_294 peakVal 't_b_294+slope' baseVal
+ t_b_295 baseVal 't_b_295+slope' peakVal
+ t_b_296 peakVal 't_b_296+slope' baseVal
+ t_b_297 baseVal 't_b_297+slope' peakVal
+ t_b_298 peakVal 't_b_298+slope' baseVal
+ t_b_299 baseVal 't_b_299+slope' peakVal
+ t_b_300 peakVal 't_b_300+slope' baseVal
+ t_b_301 baseVal 't_b_301+slope' peakVal
+ t_b_302 peakVal 't_b_302+slope' baseVal
+ t_b_303 baseVal 't_b_303+slope' peakVal
+ t_b_304 peakVal 't_b_304+slope' baseVal
+ t_b_305 baseVal 't_b_305+slope' peakVal
+ t_b_306 peakVal 't_b_306+slope' baseVal
+ t_b_307 baseVal 't_b_307+slope' peakVal
+ t_b_308 peakVal 't_b_308+slope' baseVal
+ t_b_309 baseVal 't_b_309+slope' peakVal
+ t_b_310 peakVal 't_b_310+slope' baseVal
+ t_b_311 baseVal 't_b_311+slope' peakVal
+ t_b_312 peakVal 't_b_312+slope' baseVal
+ t_b_313 baseVal 't_b_313+slope' peakVal
+ t_b_314 peakVal 't_b_314+slope' baseVal
+ t_b_315 baseVal 't_b_315+slope' peakVal
+ t_b_316 peakVal 't_b_316+slope' baseVal
+ t_b_317 baseVal 't_b_317+slope' peakVal
+ t_b_318 peakVal 't_b_318+slope' baseVal
+ t_b_319 baseVal 't_b_319+slope' peakVal
+ t_b_320 peakVal 't_b_320+slope' baseVal
+ t_b_321 baseVal 't_b_321+slope' peakVal
+ t_b_322 peakVal 't_b_322+slope' baseVal
+ t_b_323 baseVal 't_b_323+slope' peakVal
+ t_b_324 peakVal 't_b_324+slope' baseVal
+ t_b_325 baseVal 't_b_325+slope' peakVal
+ t_b_326 peakVal 't_b_326+slope' baseVal
+ t_b_327 baseVal 't_b_327+slope' peakVal
+ t_b_328 peakVal 't_b_328+slope' baseVal
+ t_b_329 baseVal 't_b_329+slope' peakVal
+ t_b_330 peakVal 't_b_330+slope' baseVal
+ t_b_331 baseVal 't_b_331+slope' peakVal
+ t_b_332 peakVal 't_b_332+slope' baseVal
+ t_b_333 baseVal 't_b_333+slope' peakVal
+ t_b_334 peakVal 't_b_334+slope' baseVal
+ t_b_335 baseVal 't_b_335+slope' peakVal
+ t_b_336 peakVal 't_b_336+slope' baseVal
+ t_b_337 baseVal 't_b_337+slope' peakVal
+ t_b_338 peakVal 't_b_338+slope' baseVal
+ t_b_339 baseVal 't_b_339+slope' peakVal
+ t_b_340 peakVal 't_b_340+slope' baseVal
+ t_b_341 baseVal 't_b_341+slope' peakVal
+ t_b_342 peakVal 't_b_342+slope' baseVal
+ t_b_343 baseVal 't_b_343+slope' peakVal
+ t_b_344 peakVal 't_b_344+slope' baseVal
+ t_b_345 baseVal 't_b_345+slope' peakVal
+ t_b_346 peakVal 't_b_346+slope' baseVal
+ t_b_347 baseVal 't_b_347+slope' peakVal
+ t_b_348 peakVal 't_b_348+slope' baseVal
+ t_b_349 baseVal 't_b_349+slope' peakVal
+ t_b_350 peakVal 't_b_350+slope' baseVal
+ t_b_351 baseVal 't_b_351+slope' peakVal
+ t_b_352 peakVal 't_b_352+slope' baseVal
+ t_b_353 baseVal 't_b_353+slope' peakVal
+ t_b_354 peakVal 't_b_354+slope' baseVal
+ t_b_355 baseVal 't_b_355+slope' peakVal
+ t_b_356 peakVal 't_b_356+slope' baseVal
+ t_b_357 baseVal 't_b_357+slope' peakVal
+ t_b_358 peakVal 't_b_358+slope' baseVal
+ t_b_359 baseVal 't_b_359+slope' peakVal
+ t_b_360 peakVal 't_b_360+slope' baseVal
+ t_b_361 baseVal 't_b_361+slope' peakVal
+ t_b_362 peakVal 't_b_362+slope' baseVal
+ t_b_363 baseVal 't_b_363+slope' peakVal
+ t_b_364 peakVal 't_b_364+slope' baseVal
+ t_b_365 baseVal 't_b_365+slope' peakVal
+ t_b_366 peakVal 't_b_366+slope' baseVal
+ t_b_367 baseVal 't_b_367+slope' peakVal
+ t_b_368 peakVal 't_b_368+slope' baseVal
+ t_b_369 baseVal 't_b_369+slope' peakVal
+ t_b_370 peakVal 't_b_370+slope' baseVal
+ t_b_371 baseVal 't_b_371+slope' peakVal
+ t_b_372 peakVal 't_b_372+slope' baseVal
+ t_b_373 baseVal 't_b_373+slope' peakVal
+ t_b_374 peakVal 't_b_374+slope' baseVal
+ t_b_375 baseVal 't_b_375+slope' peakVal
+ t_b_376 peakVal 't_b_376+slope' baseVal
+ t_b_377 baseVal 't_b_377+slope' peakVal
+ t_b_378 peakVal 't_b_378+slope' baseVal
+ t_b_379 baseVal 't_b_379+slope' peakVal
+ t_b_380 peakVal 't_b_380+slope' baseVal
+ t_b_381 baseVal 't_b_381+slope' peakVal
+ t_b_382 peakVal 't_b_382+slope' baseVal
+ t_b_383 baseVal 't_b_383+slope' peakVal
+ t_b_384 peakVal 't_b_384+slope' baseVal
+ t_b_385 baseVal 't_b_385+slope' peakVal
+ t_b_386 peakVal 't_b_386+slope' baseVal
+ t_b_387 baseVal 't_b_387+slope' peakVal
+ t_b_388 peakVal 't_b_388+slope' baseVal
+ t_b_389 baseVal 't_b_389+slope' peakVal
+ t_b_390 peakVal 't_b_390+slope' baseVal
+ t_b_391 baseVal 't_b_391+slope' peakVal
+ t_b_392 peakVal 't_b_392+slope' baseVal
+ t_b_393 baseVal 't_b_393+slope' peakVal
+ t_b_394 peakVal 't_b_394+slope' baseVal
+ t_b_395 baseVal 't_b_395+slope' peakVal
+ t_b_396 peakVal 't_b_396+slope' baseVal
+ t_b_397 baseVal 't_b_397+slope' peakVal
+ t_b_398 peakVal 't_b_398+slope' baseVal
+ t_b_399 baseVal 't_b_399+slope' peakVal
+ t_b_400 peakVal 't_b_400+slope' baseVal
+ t_b_401 baseVal 't_b_401+slope' peakVal
+ t_b_402 peakVal 't_b_402+slope' baseVal
+ t_b_403 baseVal 't_b_403+slope' peakVal
+ t_b_404 peakVal 't_b_404+slope' baseVal
+ t_b_405 baseVal 't_b_405+slope' peakVal
+ t_b_406 peakVal 't_b_406+slope' baseVal
+ t_b_407 baseVal 't_b_407+slope' peakVal
+ t_b_408 peakVal 't_b_408+slope' baseVal
+ t_b_409 baseVal 't_b_409+slope' peakVal
+ t_b_410 peakVal 't_b_410+slope' baseVal
+ t_b_411 baseVal 't_b_411+slope' peakVal
+ t_b_412 peakVal 't_b_412+slope' baseVal
+ t_b_413 baseVal 't_b_413+slope' peakVal
+ t_b_414 peakVal 't_b_414+slope' baseVal
+ t_b_415 baseVal 't_b_415+slope' peakVal
+ t_b_416 peakVal 't_b_416+slope' baseVal
+ t_b_417 baseVal 't_b_417+slope' peakVal
+ t_b_418 peakVal 't_b_418+slope' baseVal
+ t_b_419 baseVal 't_b_419+slope' peakVal
+ t_b_420 peakVal 't_b_420+slope' baseVal
+ t_b_421 baseVal 't_b_421+slope' peakVal
+ t_b_422 peakVal 't_b_422+slope' baseVal
+ t_b_423 baseVal 't_b_423+slope' peakVal
+ t_b_424 peakVal 't_b_424+slope' baseVal
+ t_b_425 baseVal 't_b_425+slope' peakVal
+ t_b_426 peakVal 't_b_426+slope' baseVal
+ t_b_427 baseVal 't_b_427+slope' peakVal
+ t_b_428 peakVal 't_b_428+slope' baseVal
+ t_b_429 baseVal 't_b_429+slope' peakVal
+ t_b_430 peakVal 't_b_430+slope' baseVal
+ t_b_431 baseVal 't_b_431+slope' peakVal
+ t_b_432 peakVal 't_b_432+slope' baseVal
+ t_b_433 baseVal 't_b_433+slope' peakVal
+ t_b_434 peakVal 't_b_434+slope' baseVal
+ t_b_435 baseVal 't_b_435+slope' peakVal
+ t_b_436 peakVal 't_b_436+slope' baseVal
+ t_b_437 baseVal 't_b_437+slope' peakVal
+ t_b_438 peakVal 't_b_438+slope' baseVal
+ t_b_439 baseVal 't_b_439+slope' peakVal
+ t_b_440 peakVal 't_b_440+slope' baseVal
+ t_b_441 baseVal 't_b_441+slope' peakVal
+ t_b_442 peakVal 't_b_442+slope' baseVal
+ t_b_443 baseVal 't_b_443+slope' peakVal
+ t_b_444 peakVal 't_b_444+slope' baseVal
+ t_b_445 baseVal 't_b_445+slope' peakVal
+ t_b_446 peakVal 't_b_446+slope' baseVal
+ t_b_447 baseVal 't_b_447+slope' peakVal
+ t_b_448 peakVal 't_b_448+slope' baseVal
+ t_b_449 baseVal 't_b_449+slope' peakVal
+ t_b_450 peakVal 't_b_450+slope' baseVal
+ t_b_451 baseVal 't_b_451+slope' peakVal
+ t_b_452 peakVal 't_b_452+slope' baseVal
+ t_b_453 baseVal 't_b_453+slope' peakVal
+ t_b_454 peakVal 't_b_454+slope' baseVal
+ t_b_455 baseVal 't_b_455+slope' peakVal
+ t_b_456 peakVal 't_b_456+slope' baseVal
+ t_b_457 baseVal 't_b_457+slope' peakVal
+ t_b_458 peakVal 't_b_458+slope' baseVal
+ t_b_459 baseVal 't_b_459+slope' peakVal
+ t_b_460 peakVal 't_b_460+slope' baseVal
+ t_b_461 baseVal 't_b_461+slope' peakVal
+ t_b_462 peakVal 't_b_462+slope' baseVal
+ t_b_463 baseVal 't_b_463+slope' peakVal
+ t_b_464 peakVal 't_b_464+slope' baseVal
+ t_b_465 baseVal 't_b_465+slope' peakVal
+ t_b_466 peakVal 't_b_466+slope' baseVal
+ t_b_467 baseVal 't_b_467+slope' peakVal
+ t_b_468 peakVal 't_b_468+slope' baseVal
+ t_b_469 baseVal 't_b_469+slope' peakVal
+ t_b_470 peakVal 't_b_470+slope' baseVal
+ t_b_471 baseVal 't_b_471+slope' peakVal
+ t_b_472 peakVal 't_b_472+slope' baseVal
+ t_b_473 baseVal 't_b_473+slope' peakVal
+ t_b_474 peakVal 't_b_474+slope' baseVal
+ t_b_475 baseVal 't_b_475+slope' peakVal
+ t_b_476 peakVal 't_b_476+slope' baseVal
+ t_b_477 baseVal 't_b_477+slope' peakVal
+ t_b_478 peakVal 't_b_478+slope' baseVal
+ t_b_479 baseVal 't_b_479+slope' peakVal
+ t_b_480 peakVal 't_b_480+slope' baseVal
+ t_b_481 baseVal 't_b_481+slope' peakVal
+ t_b_482 peakVal 't_b_482+slope' baseVal
+ t_b_483 baseVal 't_b_483+slope' peakVal
+ t_b_484 peakVal 't_b_484+slope' baseVal
+ t_b_485 baseVal 't_b_485+slope' peakVal
+ t_b_486 peakVal 't_b_486+slope' baseVal
+ t_b_487 baseVal 't_b_487+slope' peakVal
+ t_b_488 peakVal 't_b_488+slope' baseVal
+ t_b_489 baseVal 't_b_489+slope' peakVal
+ t_b_490 peakVal 't_b_490+slope' baseVal
+ t_b_491 baseVal 't_b_491+slope' peakVal
+ t_b_492 peakVal 't_b_492+slope' baseVal
+ t_b_493 baseVal 't_b_493+slope' peakVal
+ t_b_494 peakVal 't_b_494+slope' baseVal
+ t_b_495 baseVal 't_b_495+slope' peakVal
+ t_b_496 peakVal 't_b_496+slope' baseVal
+ t_b_497 baseVal 't_b_497+slope' peakVal
+ t_b_498 peakVal 't_b_498+slope' baseVal
+ t_b_499 baseVal 't_b_499+slope' peakVal
+ t_b_500 peakVal 't_b_500+slope' baseVal
+ t_b_501 baseVal 't_b_501+slope' peakVal
+ t_b_502 peakVal 't_b_502+slope' baseVal
+ t_b_503 baseVal 't_b_503+slope' peakVal
+ t_b_504 peakVal 't_b_504+slope' baseVal
+ t_b_505 baseVal 't_b_505+slope' peakVal
+ t_b_506 peakVal 't_b_506+slope' baseVal
+ t_b_507 baseVal 't_b_507+slope' peakVal
+ t_b_508 peakVal 't_b_508+slope' baseVal
+ t_b_509 baseVal 't_b_509+slope' peakVal
+ t_b_510 peakVal 't_b_510+slope' baseVal
+ t_b_511 baseVal 't_b_511+slope' peakVal
+ t_b_512 peakVal 't_b_512+slope' baseVal
+ t_b_513 baseVal 't_b_513+slope' peakVal
+ t_b_514 peakVal 't_b_514+slope' baseVal
+ t_b_515 baseVal 't_b_515+slope' peakVal
+ t_b_516 peakVal 't_b_516+slope' baseVal
+ t_b_517 baseVal 't_b_517+slope' peakVal
+ t_b_518 peakVal 't_b_518+slope' baseVal
+ t_b_519 baseVal 't_b_519+slope' peakVal
+ t_b_520 peakVal 't_b_520+slope' baseVal
+ t_b_521 baseVal 't_b_521+slope' peakVal
+ t_b_522 peakVal 't_b_522+slope' baseVal
+ t_b_523 baseVal 't_b_523+slope' peakVal
+ t_b_524 peakVal 't_b_524+slope' baseVal
+ t_b_525 baseVal 't_b_525+slope' peakVal
+ t_b_526 peakVal 't_b_526+slope' baseVal
+ t_b_527 baseVal 't_b_527+slope' peakVal
+ t_b_528 peakVal 't_b_528+slope' baseVal
+ t_b_529 baseVal 't_b_529+slope' peakVal
+ t_b_530 peakVal 't_b_530+slope' baseVal
+ t_b_531 baseVal 't_b_531+slope' peakVal
+ t_b_532 peakVal 't_b_532+slope' baseVal
+ t_b_533 baseVal 't_b_533+slope' peakVal
+ t_b_534 peakVal 't_b_534+slope' baseVal
+ t_b_535 baseVal 't_b_535+slope' peakVal
+ t_b_536 peakVal 't_b_536+slope' baseVal
+ t_b_537 baseVal 't_b_537+slope' peakVal
+ t_b_538 peakVal 't_b_538+slope' baseVal
+ t_b_539 baseVal 't_b_539+slope' peakVal
+ t_b_540 peakVal 't_b_540+slope' baseVal
+ t_b_541 baseVal 't_b_541+slope' peakVal
+ t_b_542 peakVal 't_b_542+slope' baseVal
+ t_b_543 baseVal 't_b_543+slope' peakVal
+ t_b_544 peakVal 't_b_544+slope' baseVal
+ t_b_545 baseVal 't_b_545+slope' peakVal
+ t_b_546 peakVal 't_b_546+slope' baseVal
+ t_b_547 baseVal 't_b_547+slope' peakVal
+ t_b_548 peakVal 't_b_548+slope' baseVal
+ t_b_549 baseVal 't_b_549+slope' peakVal
+ t_b_550 peakVal 't_b_550+slope' baseVal
+ t_b_551 baseVal 't_b_551+slope' peakVal
+ t_b_552 peakVal 't_b_552+slope' baseVal
+ t_b_553 baseVal 't_b_553+slope' peakVal
+ t_b_554 peakVal 't_b_554+slope' baseVal
+ t_b_555 baseVal 't_b_555+slope' peakVal
+ t_b_556 peakVal 't_b_556+slope' baseVal
+ t_b_557 baseVal 't_b_557+slope' peakVal
+ t_b_558 peakVal 't_b_558+slope' baseVal
+ t_b_559 baseVal 't_b_559+slope' peakVal
+ t_b_560 peakVal 't_b_560+slope' baseVal
+ t_b_561 baseVal 't_b_561+slope' peakVal
+ t_b_562 peakVal 't_b_562+slope' baseVal
+ t_b_563 baseVal 't_b_563+slope' peakVal
+ t_b_564 peakVal 't_b_564+slope' baseVal
+ t_b_565 baseVal 't_b_565+slope' peakVal
+ t_b_566 peakVal 't_b_566+slope' baseVal
+ t_b_567 baseVal 't_b_567+slope' peakVal
+ t_b_568 peakVal 't_b_568+slope' baseVal
+ t_b_569 baseVal 't_b_569+slope' peakVal
+ t_b_570 peakVal 't_b_570+slope' baseVal
+ t_b_571 baseVal 't_b_571+slope' peakVal
+ t_b_572 peakVal 't_b_572+slope' baseVal
+ t_b_573 baseVal 't_b_573+slope' peakVal
+ t_b_574 peakVal 't_b_574+slope' baseVal
+ t_b_575 baseVal 't_b_575+slope' peakVal
+ t_b_576 peakVal 't_b_576+slope' baseVal
+ t_b_577 baseVal 't_b_577+slope' peakVal
+ t_b_578 peakVal 't_b_578+slope' baseVal
+ t_b_579 baseVal 't_b_579+slope' peakVal
+ t_b_580 peakVal 't_b_580+slope' baseVal
+ t_b_581 baseVal 't_b_581+slope' peakVal
+ t_b_582 peakVal 't_b_582+slope' baseVal
+ t_b_583 baseVal 't_b_583+slope' peakVal
+ t_b_584 peakVal 't_b_584+slope' baseVal
+ t_b_585 baseVal 't_b_585+slope' peakVal
+ t_b_586 peakVal 't_b_586+slope' baseVal
+ t_b_587 baseVal 't_b_587+slope' peakVal
+ t_b_588 peakVal 't_b_588+slope' baseVal
+ t_b_589 baseVal 't_b_589+slope' peakVal
+ t_b_590 peakVal 't_b_590+slope' baseVal
+ t_b_591 baseVal 't_b_591+slope' peakVal
+ t_b_592 peakVal 't_b_592+slope' baseVal
+ t_b_593 baseVal 't_b_593+slope' peakVal
+ t_b_594 peakVal 't_b_594+slope' baseVal
+ t_b_595 baseVal 't_b_595+slope' peakVal
+ t_b_596 peakVal 't_b_596+slope' baseVal
+ t_b_597 baseVal 't_b_597+slope' peakVal
+ t_b_598 peakVal 't_b_598+slope' baseVal
+ t_b_599 baseVal 't_b_599+slope' peakVal
+ t_b_600 peakVal 't_b_600+slope' baseVal
+ t_b_601 baseVal 't_b_601+slope' peakVal
+ t_b_602 peakVal 't_b_602+slope' baseVal
+ t_b_603 baseVal 't_b_603+slope' peakVal
+ t_b_604 peakVal 't_b_604+slope' baseVal
+ t_b_605 baseVal 't_b_605+slope' peakVal
+ t_b_606 peakVal 't_b_606+slope' baseVal
+ t_b_607 baseVal 't_b_607+slope' peakVal
+ t_b_608 peakVal 't_b_608+slope' baseVal
+ t_b_609 baseVal 't_b_609+slope' peakVal
+ t_b_610 peakVal 't_b_610+slope' baseVal
+ t_b_611 baseVal 't_b_611+slope' peakVal
+ t_b_612 peakVal 't_b_612+slope' baseVal
+ t_b_613 baseVal 't_b_613+slope' peakVal
+ t_b_614 peakVal 't_b_614+slope' baseVal
+ t_b_615 baseVal 't_b_615+slope' peakVal
+ t_b_616 peakVal 't_b_616+slope' baseVal
+ t_b_617 baseVal 't_b_617+slope' peakVal
+ t_b_618 peakVal 't_b_618+slope' baseVal
+ t_b_619 baseVal 't_b_619+slope' peakVal
+ t_b_620 peakVal 't_b_620+slope' baseVal
+ t_b_621 baseVal 't_b_621+slope' peakVal
+ t_b_622 peakVal 't_b_622+slope' baseVal
+ t_b_623 baseVal 't_b_623+slope' peakVal
+ t_b_624 peakVal 't_b_624+slope' baseVal
+ t_b_625 baseVal 't_b_625+slope' peakVal
+ t_b_626 peakVal 't_b_626+slope' baseVal
+ t_b_627 baseVal 't_b_627+slope' peakVal
+ t_b_628 peakVal 't_b_628+slope' baseVal
+ t_b_629 baseVal 't_b_629+slope' peakVal
+ t_b_630 peakVal 't_b_630+slope' baseVal
+ t_b_631 baseVal 't_b_631+slope' peakVal
+ t_b_632 peakVal 't_b_632+slope' baseVal
+ t_b_633 baseVal 't_b_633+slope' peakVal
+ t_b_634 peakVal 't_b_634+slope' baseVal
+ t_b_635 baseVal 't_b_635+slope' peakVal
+ t_b_636 peakVal 't_b_636+slope' baseVal
+ t_b_637 baseVal 't_b_637+slope' peakVal
+ t_b_638 peakVal 't_b_638+slope' baseVal
+ t_b_639 baseVal 't_b_639+slope' peakVal
+ t_b_640 peakVal 't_b_640+slope' baseVal
+ t_b_641 baseVal 't_b_641+slope' peakVal
+ t_b_642 peakVal 't_b_642+slope' baseVal
+ t_b_643 baseVal 't_b_643+slope' peakVal
+ t_b_644 peakVal 't_b_644+slope' baseVal
+ t_b_645 baseVal 't_b_645+slope' peakVal
+ t_b_646 peakVal 't_b_646+slope' baseVal
+ t_b_647 baseVal 't_b_647+slope' peakVal
+ t_b_648 peakVal 't_b_648+slope' baseVal
+ t_b_649 baseVal 't_b_649+slope' peakVal
+ t_b_650 peakVal 't_b_650+slope' baseVal
+ t_b_651 baseVal 't_b_651+slope' peakVal
+ t_b_652 peakVal 't_b_652+slope' baseVal
+ t_b_653 baseVal 't_b_653+slope' peakVal
+ t_b_654 peakVal 't_b_654+slope' baseVal
+ t_b_655 baseVal 't_b_655+slope' peakVal
+ t_b_656 peakVal 't_b_656+slope' baseVal
+ t_b_657 baseVal 't_b_657+slope' peakVal
+ t_b_658 peakVal 't_b_658+slope' baseVal
+ t_b_659 baseVal 't_b_659+slope' peakVal
+ t_b_660 peakVal 't_b_660+slope' baseVal
+ t_b_661 baseVal 't_b_661+slope' peakVal
+ t_b_662 peakVal 't_b_662+slope' baseVal
+ t_b_663 baseVal 't_b_663+slope' peakVal
+ t_b_664 peakVal 't_b_664+slope' baseVal
+ t_b_665 baseVal 't_b_665+slope' peakVal
+ t_b_666 peakVal 't_b_666+slope' baseVal
+ t_b_667 baseVal 't_b_667+slope' peakVal
+ t_b_668 peakVal 't_b_668+slope' baseVal
+ t_b_669 baseVal 't_b_669+slope' peakVal
+ t_b_670 peakVal 't_b_670+slope' baseVal
+ t_b_671 baseVal 't_b_671+slope' peakVal
+ t_b_672 peakVal 't_b_672+slope' baseVal
+ t_b_673 baseVal 't_b_673+slope' peakVal
+ t_b_674 peakVal 't_b_674+slope' baseVal
+ t_b_675 baseVal 't_b_675+slope' peakVal
+ t_b_676 peakVal 't_b_676+slope' baseVal
+ t_b_677 baseVal 't_b_677+slope' peakVal
+ t_b_678 peakVal 't_b_678+slope' baseVal
+ t_b_679 baseVal 't_b_679+slope' peakVal
+ t_b_680 peakVal 't_b_680+slope' baseVal
+ t_b_681 baseVal 't_b_681+slope' peakVal
+ t_b_682 peakVal 't_b_682+slope' baseVal
+ t_b_683 baseVal 't_b_683+slope' peakVal
+ t_b_684 peakVal 't_b_684+slope' baseVal
+ t_b_685 baseVal 't_b_685+slope' peakVal
+ t_b_686 peakVal 't_b_686+slope' baseVal
+ t_b_687 baseVal 't_b_687+slope' peakVal
+ t_b_688 peakVal 't_b_688+slope' baseVal
+ t_b_689 baseVal 't_b_689+slope' peakVal
+ t_b_690 peakVal 't_b_690+slope' baseVal
+ t_b_691 baseVal 't_b_691+slope' peakVal
+ t_b_692 peakVal 't_b_692+slope' baseVal
+ t_b_693 baseVal 't_b_693+slope' peakVal
+ t_b_694 peakVal 't_b_694+slope' baseVal
+ t_b_695 baseVal 't_b_695+slope' peakVal
+ t_b_696 peakVal 't_b_696+slope' baseVal
+ t_b_697 baseVal 't_b_697+slope' peakVal
+ t_b_698 peakVal 't_b_698+slope' baseVal
+ t_b_699 baseVal 't_b_699+slope' peakVal
+ t_b_700 peakVal 't_b_700+slope' baseVal
+ t_b_701 baseVal 't_b_701+slope' peakVal
+ t_b_702 peakVal 't_b_702+slope' baseVal
+ t_b_703 baseVal 't_b_703+slope' peakVal
+ t_b_704 peakVal 't_b_704+slope' baseVal
+ t_b_705 baseVal 't_b_705+slope' peakVal
+ t_b_706 peakVal 't_b_706+slope' baseVal
+ t_b_707 baseVal 't_b_707+slope' peakVal
+ t_b_708 peakVal 't_b_708+slope' baseVal
+ t_b_709 baseVal 't_b_709+slope' peakVal
+ t_b_710 peakVal 't_b_710+slope' baseVal
+ t_b_711 baseVal 't_b_711+slope' peakVal
+ t_b_712 peakVal 't_b_712+slope' baseVal
+ t_b_713 baseVal 't_b_713+slope' peakVal
+ t_b_714 peakVal 't_b_714+slope' baseVal
+ t_b_715 baseVal 't_b_715+slope' peakVal
+ t_b_716 peakVal 't_b_716+slope' baseVal
+ t_b_717 baseVal 't_b_717+slope' peakVal
+ t_b_718 peakVal 't_b_718+slope' baseVal
+ t_b_719 baseVal 't_b_719+slope' peakVal
+ t_b_720 peakVal 't_b_720+slope' baseVal
+ t_b_721 baseVal 't_b_721+slope' peakVal
+ t_b_722 peakVal 't_b_722+slope' baseVal
+ t_b_723 baseVal 't_b_723+slope' peakVal
+ t_b_724 peakVal 't_b_724+slope' baseVal
+ t_b_725 baseVal 't_b_725+slope' peakVal
+ t_b_726 peakVal 't_b_726+slope' baseVal
+ t_b_727 baseVal 't_b_727+slope' peakVal
+ t_b_728 peakVal 't_b_728+slope' baseVal
+ t_b_729 baseVal 't_b_729+slope' peakVal
+ t_b_730 peakVal 't_b_730+slope' baseVal
+ t_b_731 baseVal 't_b_731+slope' peakVal
+ t_b_732 peakVal 't_b_732+slope' baseVal
+ t_b_733 baseVal 't_b_733+slope' peakVal
+ t_b_734 peakVal 't_b_734+slope' baseVal
+ t_b_735 baseVal 't_b_735+slope' peakVal
+ t_b_736 peakVal 't_b_736+slope' baseVal
+ t_b_737 baseVal 't_b_737+slope' peakVal
+ t_b_738 peakVal 't_b_738+slope' baseVal
+ t_b_739 baseVal 't_b_739+slope' peakVal
+ t_b_740 peakVal 't_b_740+slope' baseVal
+ t_b_741 baseVal 't_b_741+slope' peakVal
+ t_b_742 peakVal 't_b_742+slope' baseVal
+ t_b_743 baseVal 't_b_743+slope' peakVal
+ t_b_744 peakVal 't_b_744+slope' baseVal
+ t_b_745 baseVal 't_b_745+slope' peakVal
+ t_b_746 peakVal 't_b_746+slope' baseVal
+ t_b_747 baseVal 't_b_747+slope' peakVal
+ t_b_748 peakVal 't_b_748+slope' baseVal
+ t_b_749 baseVal 't_b_749+slope' peakVal
+ t_b_750 peakVal 't_b_750+slope' baseVal
+ t_b_751 baseVal 't_b_751+slope' peakVal
+ t_b_752 peakVal 't_b_752+slope' baseVal
+ t_b_753 baseVal 't_b_753+slope' peakVal
+ t_b_754 peakVal 't_b_754+slope' baseVal
+ t_b_755 baseVal 't_b_755+slope' peakVal
+ t_b_756 peakVal 't_b_756+slope' baseVal
+ t_b_757 baseVal 't_b_757+slope' peakVal
+ t_b_758 peakVal 't_b_758+slope' baseVal
+ t_b_759 baseVal 't_b_759+slope' peakVal
+ t_b_760 peakVal 't_b_760+slope' baseVal
+ t_b_761 baseVal 't_b_761+slope' peakVal
+ t_b_762 peakVal 't_b_762+slope' baseVal
+ t_b_763 baseVal 't_b_763+slope' peakVal
+ t_b_764 peakVal 't_b_764+slope' baseVal
+ t_b_765 baseVal 't_b_765+slope' peakVal
+ t_b_766 peakVal 't_b_766+slope' baseVal
+ t_b_767 baseVal 't_b_767+slope' peakVal
+ t_b_768 peakVal 't_b_768+slope' baseVal
+ t_b_769 baseVal 't_b_769+slope' peakVal
+ t_b_770 peakVal 't_b_770+slope' baseVal
+ t_b_771 baseVal 't_b_771+slope' peakVal
+ t_b_772 peakVal 't_b_772+slope' baseVal
+ t_b_773 baseVal 't_b_773+slope' peakVal
+ t_b_774 peakVal 't_b_774+slope' baseVal
+ t_b_775 baseVal 't_b_775+slope' peakVal
+ t_b_776 peakVal 't_b_776+slope' baseVal
+ t_b_777 baseVal 't_b_777+slope' peakVal
+ t_b_778 peakVal 't_b_778+slope' baseVal
+ t_b_779 baseVal 't_b_779+slope' peakVal
+ t_b_780 peakVal 't_b_780+slope' baseVal
+ t_b_781 baseVal 't_b_781+slope' peakVal
+ t_b_782 peakVal 't_b_782+slope' baseVal
+ t_b_783 baseVal 't_b_783+slope' peakVal
+ t_b_784 peakVal 't_b_784+slope' baseVal
+ t_b_785 baseVal 't_b_785+slope' peakVal
+ t_b_786 peakVal 't_b_786+slope' baseVal
+ t_b_787 baseVal 't_b_787+slope' peakVal
+ t_b_788 peakVal 't_b_788+slope' baseVal
+ t_b_789 baseVal 't_b_789+slope' peakVal
+ t_b_790 peakVal 't_b_790+slope' baseVal
+ t_b_791 baseVal 't_b_791+slope' peakVal
+ t_b_792 peakVal 't_b_792+slope' baseVal
+ t_b_793 baseVal 't_b_793+slope' peakVal
+ t_b_794 peakVal 't_b_794+slope' baseVal
+ t_b_795 baseVal 't_b_795+slope' peakVal
+ t_b_796 peakVal 't_b_796+slope' baseVal
+ t_b_797 baseVal 't_b_797+slope' peakVal
+ t_b_798 peakVal 't_b_798+slope' baseVal
+ t_b_799 baseVal 't_b_799+slope' peakVal

*circuit

XBUFFER_A Input_A A VDD VDD GND GND BUF_X8
XBUFFER_B Input_B B VDD VDD GND GND BUF_X8
XCGATE A B Z VDD VDD GND GND CGATE
XBUFFER_Z Z Output VDD VDD GND GND BUF_X8
C_TERM Output GND 0.0779pF

.PROBE TRAN V(A) V(B) V(Z)
.TRAN 0.1ps tend
.END
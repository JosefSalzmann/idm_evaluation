* circuit: nor inv chain
simulator lang=spice

*.PARAM pw=<sed>pw<sed>as
.PARAM supp=0.8V slope=0.1fs
.PARAM t_init0=0.1ns t_init1=0.174ns
.PARAM baseVal=0V peakVal=0.8V tend=1.0ns


.LIB /home/s11777724/involution_tool_library_files/backend/spice/fet.inc CMG

* main circuit
.INCLUDE /home/s11777724/involution_tool_library_files/backend/spice/cell/INV_X1.sp

**** SPECTRE Back Annotation
.option spef='../place_and_route/generic_parasitics.spef'
****

.TEMP 25
.OPTION
+ INGOLD=2
+ PARHIER=LOCAL
*+ POST=CSDF
+ PROBE
+ BRIEF
+ ACCURATE
+ ABSVAR=0.0001
+ DVDT=2
+ RELTOL=1e-11
*+ DELMAX=100fs
+ dc_pivot_check=yes

* vdd
VDD VDD GND 0.8v

VIN myin GND PWL 0ns baseVal t_init0 baseVal 't_init0+slope' peakVal t_init1 peakVal 't_init1+slope' baseVal

* circuit under test
XINV0 myin STAGE0 VDD VDD GND GND INV_X1
XINV1 STAGE0 STAGE1 VDD VDD GND GND INV_X1
XINV2 STAGE1 STAGE2 VDD VDD GND GND INV_X1
XINV3 STAGE2 STAGE3 VDD VDD GND GND INV_X1
XINV4 STAGE3 STAGE4 VDD VDD GND GND INV_X1
XINV5 STAGE4 STAGE5 VDD VDD GND GND INV_X1
XINV6 STAGE5 STAGE6 VDD VDD GND GND INV_X1
XINV7 STAGE6 STAGE7 VDD VDD GND GND INV_X1
XINV8 STAGE7 STAGE8 VDD VDD GND GND INV_X1
XINV9 STAGE8 STAGE9 VDD VDD GND GND INV_X1
XINV10 STAGE9 STAGE10 VDD VDD GND GND INV_X1
XINV11 STAGE10 STAGE11 VDD VDD GND GND INV_X1
XINV12 STAGE11 STAGE12 VDD VDD GND GND INV_X1
XINV13 STAGE12 STAGE13 VDD VDD GND GND INV_X1
XINV14 STAGE13 STAGE14 VDD VDD GND GND INV_X1
XINV15 STAGE14 STAGE15 VDD VDD GND GND INV_X1
XINV16 STAGE15 STAGE16 VDD VDD GND GND INV_X1
XINV17 STAGE16 STAGE17 VDD VDD GND GND INV_X1
XINV18 STAGE17 STAGE18 VDD VDD GND GND INV_X1
XINV19 STAGE18 STAGE19 VDD VDD GND GND INV_X1
XINV20 STAGE19 STAGE20 VDD VDD GND GND INV_X1
XINV21 STAGE20 STAGE21 VDD VDD GND GND INV_X1
XINV22 STAGE21 STAGE22 VDD VDD GND GND INV_X1
XINV23 STAGE22 STAGE23 VDD VDD GND GND INV_X1
XINV24 STAGE23 STAGE24 VDD VDD GND GND INV_X1
XINV25 STAGE24 O_C_TERM VDD VDD GND GND INV_X1
C_TERM O_C_TERM GND 0.0779pF

.PROBE TRAN V(myin) V(STAGE0) V(STAGE1) V(STAGE2) V(STAGE3) V(STAGE4)
+ V(STAGE5) V(STAGE6) V(STAGE7) V(STAGE8) V(STAGE9) V(STAGE10)
+ V(STAGE11) V(STAGE12) V(STAGE13) V(STAGE14) V(STAGE15)
+ V(STAGE16) V(STAGE17) V(STAGE18) V(STAGE19) V(STAGE20)
+ V(STAGE21) V(STAGE22) V(STAGE23) V(STAGE24) V(O_C_TERM)
.TRAN 0.1ps tend
.END

* circuit: inv chain
simulator lang=spice

*.PARAM pw=<sed>pw<sed>as
.PARAM supp=0.8V slope=0.1fs
.PARAM t_init0=0.1ns t_init1=0.174ns
.PARAM baseVal=0V peakVal=0.8V tend=1.0ns


.LIB /home/s11777724/involution_tool_library_files/backend/spice/fet.inc CMG

* main circuit
.INCLUDE /home/s11777724/involution_tool_library_files/backend/spice/cell/INV_X1.sp

**** SPECTRE Back Annotation
.option spef='../place_and_route/generic_parasitics.spef'
****

.TEMP 25
.OPTION
+ INGOLD=2
+ PARHIER=LOCAL
*+ POST=CSDF
+ PROBE
+ BRIEF
+ ACCURATE
+ ABSVAR=0.0001
+ DVDT=2
+ RELTOL=1e-11
*+ DELMAX=100fs
+ dc_pivot_check=yes

* vdd
VDD VDD GND 0.8v

VIN myin GND PWL 0ns baseVal t_init0 baseVal 't_init0+slope' peakVal t_init1 peakVal 't_init1+slope' baseVal

* circuit under test
XINV0 myin STAGE0 VDD VDD GND GND INV_X1
XINV1 STAGE0 STAGE1 VDD VDD GND GND INV_X1
XINV2 STAGE1 STAGE2 VDD VDD GND GND INV_X1
XINV3 STAGE2 STAGE3 VDD VDD GND GND INV_X1
XINV4 STAGE3 STAGE4 VDD VDD GND GND INV_X1
XINV5 STAGE4 STAGE5 VDD VDD GND GND INV_X1
XINV6 STAGE5 STAGE6 VDD VDD GND GND INV_X1
XINV7 STAGE6 STAGE7 VDD VDD GND GND INV_X1
XINV8 STAGE7 STAGE8 VDD VDD GND GND INV_X1
XINV9 STAGE8 STAGE9 VDD VDD GND GND INV_X1
XINV10 STAGE9 STAGE10 VDD VDD GND GND INV_X1
XINV11 STAGE10 STAGE11 VDD VDD GND GND INV_X1
XINV12 STAGE11 STAGE12 VDD VDD GND GND INV_X1
XINV13 STAGE12 STAGE13 VDD VDD GND GND INV_X1
XINV14 STAGE13 STAGE14 VDD VDD GND GND INV_X1
XINV15 STAGE14 STAGE15 VDD VDD GND GND INV_X1
XINV16 STAGE15 STAGE16 VDD VDD GND GND INV_X1
XINV17 STAGE16 STAGE17 VDD VDD GND GND INV_X1
XINV18 STAGE17 STAGE18 VDD VDD GND GND INV_X1
XINV19 STAGE18 STAGE19 VDD VDD GND GND INV_X1
XINV20 STAGE19 STAGE20 VDD VDD GND GND INV_X1
XINV21 STAGE20 STAGE21 VDD VDD GND GND INV_X1
XINV22 STAGE21 STAGE22 VDD VDD GND GND INV_X1
XINV23 STAGE22 STAGE23 VDD VDD GND GND INV_X1
XINV24 STAGE23 STAGE24 VDD VDD GND GND INV_X1
XINV25 STAGE24 STAGE25 VDD VDD GND GND INV_X1
XINV26 STAGE25 STAGE26 VDD VDD GND GND INV_X1
XINV27 STAGE26 STAGE27 VDD VDD GND GND INV_X1
XINV28 STAGE27 STAGE28 VDD VDD GND GND INV_X1
XINV29 STAGE28 STAGE29 VDD VDD GND GND INV_X1
XINV30 STAGE29 STAGE30 VDD VDD GND GND INV_X1
XINV31 STAGE30 STAGE31 VDD VDD GND GND INV_X1
XINV32 STAGE31 STAGE32 VDD VDD GND GND INV_X1
XINV33 STAGE32 STAGE33 VDD VDD GND GND INV_X1
XINV34 STAGE33 STAGE34 VDD VDD GND GND INV_X1
XINV35 STAGE34 STAGE35 VDD VDD GND GND INV_X1
XINV36 STAGE35 STAGE36 VDD VDD GND GND INV_X1
XINV37 STAGE36 STAGE37 VDD VDD GND GND INV_X1
XINV38 STAGE37 STAGE38 VDD VDD GND GND INV_X1
XINV39 STAGE38 STAGE39 VDD VDD GND GND INV_X1
XINV40 STAGE39 STAGE40 VDD VDD GND GND INV_X1
XINV41 STAGE40 STAGE41 VDD VDD GND GND INV_X1
XINV42 STAGE41 STAGE42 VDD VDD GND GND INV_X1
XINV43 STAGE42 STAGE43 VDD VDD GND GND INV_X1
XINV44 STAGE43 STAGE44 VDD VDD GND GND INV_X1
XINV45 STAGE44 STAGE45 VDD VDD GND GND INV_X1
XINV46 STAGE45 STAGE46 VDD VDD GND GND INV_X1
XINV47 STAGE46 STAGE47 VDD VDD GND GND INV_X1
XINV48 STAGE47 STAGE48 VDD VDD GND GND INV_X1
XINV49 STAGE48 STAGE49 VDD VDD GND GND INV_X1
XINV50 STAGE49 STAGE50 VDD VDD GND GND INV_X1
XINV51 STAGE50 STAGE51 VDD VDD GND GND INV_X1
XINV52 STAGE51 STAGE52 VDD VDD GND GND INV_X1
XINV53 STAGE52 STAGE53 VDD VDD GND GND INV_X1
XINV54 STAGE53 STAGE54 VDD VDD GND GND INV_X1
XINV55 STAGE54 STAGE55 VDD VDD GND GND INV_X1
XINV56 STAGE55 STAGE56 VDD VDD GND GND INV_X1
XINV57 STAGE56 STAGE57 VDD VDD GND GND INV_X1
XINV58 STAGE57 STAGE58 VDD VDD GND GND INV_X1
XINV59 STAGE58 STAGE59 VDD VDD GND GND INV_X1
XINV60 STAGE59 STAGE60 VDD VDD GND GND INV_X1
XINV61 STAGE60 STAGE61 VDD VDD GND GND INV_X1
XINV62 STAGE61 STAGE62 VDD VDD GND GND INV_X1
XINV63 STAGE62 STAGE63 VDD VDD GND GND INV_X1
XINV64 STAGE63 STAGE64 VDD VDD GND GND INV_X1
XINV65 STAGE64 STAGE65 VDD VDD GND GND INV_X1
XINV66 STAGE65 STAGE66 VDD VDD GND GND INV_X1
XINV67 STAGE66 STAGE67 VDD VDD GND GND INV_X1
XINV68 STAGE67 STAGE68 VDD VDD GND GND INV_X1
XINV69 STAGE68 STAGE69 VDD VDD GND GND INV_X1
XINV70 STAGE69 STAGE70 VDD VDD GND GND INV_X1
XINV71 STAGE70 STAGE71 VDD VDD GND GND INV_X1
XINV72 STAGE71 STAGE72 VDD VDD GND GND INV_X1
XINV73 STAGE72 STAGE73 VDD VDD GND GND INV_X1
XINV74 STAGE73 STAGE74 VDD VDD GND GND INV_X1
XINV75 STAGE74 STAGE75 VDD VDD GND GND INV_X1
XINV76 STAGE75 STAGE76 VDD VDD GND GND INV_X1
XINV77 STAGE76 STAGE77 VDD VDD GND GND INV_X1
XINV78 STAGE77 STAGE78 VDD VDD GND GND INV_X1
XINV79 STAGE78 STAGE79 VDD VDD GND GND INV_X1
XINV80 STAGE79 STAGE80 VDD VDD GND GND INV_X1
XINV81 STAGE80 STAGE81 VDD VDD GND GND INV_X1
XINV82 STAGE81 STAGE82 VDD VDD GND GND INV_X1
XINV83 STAGE82 STAGE83 VDD VDD GND GND INV_X1
XINV84 STAGE83 STAGE84 VDD VDD GND GND INV_X1
XINV85 STAGE84 STAGE85 VDD VDD GND GND INV_X1
XINV86 STAGE85 STAGE86 VDD VDD GND GND INV_X1
XINV87 STAGE86 STAGE87 VDD VDD GND GND INV_X1
XINV88 STAGE87 STAGE88 VDD VDD GND GND INV_X1
XINV89 STAGE88 STAGE89 VDD VDD GND GND INV_X1
XINV90 STAGE89 STAGE90 VDD VDD GND GND INV_X1
XINV91 STAGE90 STAGE91 VDD VDD GND GND INV_X1
XINV92 STAGE91 STAGE92 VDD VDD GND GND INV_X1
XINV93 STAGE92 STAGE93 VDD VDD GND GND INV_X1
XINV94 STAGE93 STAGE94 VDD VDD GND GND INV_X1
XINV95 STAGE94 STAGE95 VDD VDD GND GND INV_X1
XINV96 STAGE95 STAGE96 VDD VDD GND GND INV_X1
XINV97 STAGE96 STAGE97 VDD VDD GND GND INV_X1
XINV98 STAGE97 STAGE98 VDD VDD GND GND INV_X1
XINV99 STAGE98 STAGE99 VDD VDD GND GND INV_X1
XINV100 STAGE99 STAGE100 VDD VDD GND GND INV_X1
XINV101 STAGE100 STAGE101 VDD VDD GND GND INV_X1
XINV102 STAGE101 STAGE102 VDD VDD GND GND INV_X1
XINV103 STAGE102 STAGE103 VDD VDD GND GND INV_X1
XINV104 STAGE103 STAGE104 VDD VDD GND GND INV_X1
XINV105 STAGE104 STAGE105 VDD VDD GND GND INV_X1
XINV106 STAGE105 STAGE106 VDD VDD GND GND INV_X1
XINV107 STAGE106 STAGE107 VDD VDD GND GND INV_X1
XINV108 STAGE107 STAGE108 VDD VDD GND GND INV_X1
XINV109 STAGE108 STAGE109 VDD VDD GND GND INV_X1
XINV110 STAGE109 STAGE110 VDD VDD GND GND INV_X1
XINV111 STAGE110 STAGE111 VDD VDD GND GND INV_X1
XINV112 STAGE111 STAGE112 VDD VDD GND GND INV_X1
XINV113 STAGE112 STAGE113 VDD VDD GND GND INV_X1
XINV114 STAGE113 STAGE114 VDD VDD GND GND INV_X1
XINV115 STAGE114 STAGE115 VDD VDD GND GND INV_X1
XINV116 STAGE115 STAGE116 VDD VDD GND GND INV_X1
XINV117 STAGE116 STAGE117 VDD VDD GND GND INV_X1
XINV118 STAGE117 STAGE118 VDD VDD GND GND INV_X1
XINV119 STAGE118 myout VDD VDD GND GND INV_X1
C_TERM myout GND 0.0779pF

.PROBE TRAN V(myin) V(STAGE1) V(STAGE2) V(STAGE3) V(STAGE4) V(STAGE5) V(STAGE6) V(STAGE7) V(STAGE8) V(STAGE9) V(STAGE10) V(STAGE11) V(STAGE12) V(STAGE13) V(STAGE14) V(STAGE15) V(STAGE16) V(STAGE17) V(STAGE18) V(STAGE19) V(STAGE20) V(STAGE21) V(STAGE22) V(STAGE23) V(STAGE24) V(STAGE25) V(STAGE26) V(STAGE27) V(STAGE28) V(STAGE29) V(STAGE30) V(STAGE31) V(STAGE32) V(STAGE33) V(STAGE34) V(STAGE35) V(STAGE36) V(STAGE37) V(STAGE38) V(STAGE39) V(STAGE40) V(STAGE41) V(STAGE42) V(STAGE43) V(STAGE44) V(STAGE45) V(STAGE46) V(STAGE47) V(STAGE48) V(STAGE49) V(STAGE50) V(STAGE51) V(STAGE52) V(STAGE53) V(STAGE54) V(STAGE55) V(STAGE56) V(STAGE57) V(STAGE58) V(STAGE59) V(STAGE60) V(STAGE61) V(STAGE62) V(STAGE63) V(STAGE64) V(STAGE65) V(STAGE66) V(STAGE67) V(STAGE68) V(STAGE69) V(STAGE70) V(STAGE71) V(STAGE72) V(STAGE73) V(STAGE74) V(STAGE75) V(STAGE76) V(STAGE77) V(STAGE78) V(STAGE79) V(STAGE80) V(STAGE81) V(STAGE82) V(STAGE83) V(STAGE84) V(STAGE85) V(STAGE86) V(STAGE87) V(STAGE88) V(STAGE89) V(STAGE90) V(STAGE91) V(STAGE92) V(STAGE93) V(STAGE94) V(STAGE95) V(STAGE96) V(STAGE97) V(STAGE98) V(STAGE99) V(STAGE100) V(STAGE101) V(STAGE102) V(STAGE103) V(STAGE104) V(STAGE105) V(STAGE106) V(STAGE107) V(STAGE108) V(STAGE109) V(STAGE110) V(STAGE111) V(STAGE112) V(STAGE113) V(STAGE114) V(STAGE115)
.TRAN 0.1ps tend
.END

module c1908_NOR_template (N1_PWL,N4_PWL,N7_PWL,N10_PWL,N13_PWL,N16_PWL,N19_PWL,N22_PWL,
            N25_PWL,N28_PWL,N31_PWL,N34_PWL,N37_PWL,N40_PWL,N43_PWL,N46_PWL,N49_PWL,
            N53_PWL,N56_PWL,N60_PWL,N63_PWL,N66_PWL,N69_PWL,N72_PWL,N76_PWL,N79_PWL,
            N82_PWL,N85_PWL,N88_PWL,N91_PWL,N94_PWL,N99_PWL,N104_PWL,
            N2753_TERMINATION,N2754_TERMINATION,N2755_TERMINATION,N2756_TERMINATION,
            N2762_TERMINATION,N2767_TERMINATION,N2768_TERMINATION,N2779_TERMINATION,
            N2780_TERMINATION,N2781_TERMINATION,N2782_TERMINATION,N2783_TERMINATION,
            N2784_TERMINATION,N2785_TERMINATION,N2786_TERMINATION,N2787_TERMINATION,
            N2811_TERMINATION,N2886_TERMINATION,N2887_TERMINATION,N2888_TERMINATION,
            N2889_TERMINATION,N2890_TERMINATION,N2891_TERMINATION,N2892_TERMINATION,
            N2899_TERMINATION);



      input N1_PWL,N4_PWL,N7_PWL,N10_PWL,N13_PWL,N16_PWL,N19_PWL,N22_PWL,
            N25_PWL,N28_PWL,N31_PWL,N34_PWL,N37_PWL,N40_PWL,N43_PWL,N46_PWL,N49_PWL,
            N53_PWL,N56_PWL,N60_PWL,N63_PWL,N66_PWL,N69_PWL,N72_PWL,N76_PWL,N79_PWL,
            N82_PWL,N85_PWL,N88_PWL,N91_PWL,N94_PWL,N99_PWL,N104_PWL;

      output N2753_TERMINATION,N2754_TERMINATION,N2755_TERMINATION,N2756_TERMINATION,
            N2762_TERMINATION,N2767_TERMINATION,N2768_TERMINATION,N2779_TERMINATION,
            N2780_TERMINATION,N2781_TERMINATION,N2782_TERMINATION,N2783_TERMINATION,
            N2784_TERMINATION,N2785_TERMINATION,N2786_TERMINATION,N2787_TERMINATION,
            N2811_TERMINATION,N2886_TERMINATION,N2887_TERMINATION,N2888_TERMINATION,
            N2889_TERMINATION,N2890_TERMINATION,N2891_TERMINATION,N2892_TERMINATION,
            N2899_TERMINATION;

      wire GND = 1'b0;
      wire XNOR_1_1_N1_PULSESHAPING_OUT, XNOR_1_2_N1_PULSESHAPING_OUT, XNOR_1_3_N1_PULSESHAPING_OUT, XNOR_1_4_N1_PULSESHAPING_OUT, XNOR_1_5_N1_PULSESHAPING_OUT, XNOR_1_6_N1_PULSESHAPING_OUT;
      NOR2_X1 XNOR_1_1_N1_PULSESHAPING (.ZN (XNOR_1_1_N1_PULSESHAPING_OUT), .A1 (N1_PWL), .A2 (GND));
      NOR2_X1 XNOR_1_2_N1_PULSESHAPING (.ZN (XNOR_1_2_N1_PULSESHAPING_OUT), .A1 (XNOR_1_1_N1_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_3_N1_PULSESHAPING (.ZN (XNOR_1_3_N1_PULSESHAPING_OUT), .A1 (XNOR_1_2_N1_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_4_N1_PULSESHAPING (.ZN (XNOR_1_4_N1_PULSESHAPING_OUT), .A1 (XNOR_1_3_N1_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_5_N1_PULSESHAPING (.ZN (XNOR_1_5_N1_PULSESHAPING_OUT), .A1 (XNOR_1_4_N1_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_6_N1_PULSESHAPING (.ZN (XNOR_1_6_N1_PULSESHAPING_OUT), .A1 (XNOR_1_5_N1_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_7_N1_PULSESHAPING (.ZN (N1), .A1 (XNOR_1_6_N1_PULSESHAPING_OUT), .A2 (GND));

      wire XNOR_1_1_N4_PULSESHAPING_OUT, XNOR_1_2_N4_PULSESHAPING_OUT, XNOR_1_3_N4_PULSESHAPING_OUT, XNOR_1_4_N4_PULSESHAPING_OUT, XNOR_1_5_N4_PULSESHAPING_OUT, XNOR_1_6_N4_PULSESHAPING_OUT;
      NOR2_X1 XNOR_1_1_N4_PULSESHAPING (.ZN (XNOR_1_1_N4_PULSESHAPING_OUT), .A1 (N4_PWL), .A2 (GND));
      NOR2_X1 XNOR_1_2_N4_PULSESHAPING (.ZN (XNOR_1_2_N4_PULSESHAPING_OUT), .A1 (XNOR_1_1_N4_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_3_N4_PULSESHAPING (.ZN (XNOR_1_3_N4_PULSESHAPING_OUT), .A1 (XNOR_1_2_N4_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_4_N4_PULSESHAPING (.ZN (XNOR_1_4_N4_PULSESHAPING_OUT), .A1 (XNOR_1_3_N4_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_5_N4_PULSESHAPING (.ZN (XNOR_1_5_N4_PULSESHAPING_OUT), .A1 (XNOR_1_4_N4_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_6_N4_PULSESHAPING (.ZN (XNOR_1_6_N4_PULSESHAPING_OUT), .A1 (XNOR_1_5_N4_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_7_N4_PULSESHAPING (.ZN (N4), .A1 (XNOR_1_6_N4_PULSESHAPING_OUT), .A2 (GND));

      wire XNOR_1_1_N7_PULSESHAPING_OUT, XNOR_1_2_N7_PULSESHAPING_OUT, XNOR_1_3_N7_PULSESHAPING_OUT, XNOR_1_4_N7_PULSESHAPING_OUT, XNOR_1_5_N7_PULSESHAPING_OUT, XNOR_1_6_N7_PULSESHAPING_OUT;
      NOR2_X1 XNOR_1_1_N7_PULSESHAPING (.ZN (XNOR_1_1_N7_PULSESHAPING_OUT), .A1 (N7_PWL), .A2 (GND));
      NOR2_X1 XNOR_1_2_N7_PULSESHAPING (.ZN (XNOR_1_2_N7_PULSESHAPING_OUT), .A1 (XNOR_1_1_N7_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_3_N7_PULSESHAPING (.ZN (XNOR_1_3_N7_PULSESHAPING_OUT), .A1 (XNOR_1_2_N7_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_4_N7_PULSESHAPING (.ZN (XNOR_1_4_N7_PULSESHAPING_OUT), .A1 (XNOR_1_3_N7_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_5_N7_PULSESHAPING (.ZN (XNOR_1_5_N7_PULSESHAPING_OUT), .A1 (XNOR_1_4_N7_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_6_N7_PULSESHAPING (.ZN (XNOR_1_6_N7_PULSESHAPING_OUT), .A1 (XNOR_1_5_N7_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_7_N7_PULSESHAPING (.ZN (N7), .A1 (XNOR_1_6_N7_PULSESHAPING_OUT), .A2 (GND));

      wire XNOR_1_1_N10_PULSESHAPING_OUT, XNOR_1_2_N10_PULSESHAPING_OUT, XNOR_1_3_N10_PULSESHAPING_OUT, XNOR_1_4_N10_PULSESHAPING_OUT, XNOR_1_5_N10_PULSESHAPING_OUT, XNOR_1_6_N10_PULSESHAPING_OUT;
      NOR2_X1 XNOR_1_1_N10_PULSESHAPING (.ZN (XNOR_1_1_N10_PULSESHAPING_OUT), .A1 (N10_PWL), .A2 (GND));
      NOR2_X1 XNOR_1_2_N10_PULSESHAPING (.ZN (XNOR_1_2_N10_PULSESHAPING_OUT), .A1 (XNOR_1_1_N10_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_3_N10_PULSESHAPING (.ZN (XNOR_1_3_N10_PULSESHAPING_OUT), .A1 (XNOR_1_2_N10_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_4_N10_PULSESHAPING (.ZN (XNOR_1_4_N10_PULSESHAPING_OUT), .A1 (XNOR_1_3_N10_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_5_N10_PULSESHAPING (.ZN (XNOR_1_5_N10_PULSESHAPING_OUT), .A1 (XNOR_1_4_N10_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_6_N10_PULSESHAPING (.ZN (XNOR_1_6_N10_PULSESHAPING_OUT), .A1 (XNOR_1_5_N10_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_7_N10_PULSESHAPING (.ZN (N10), .A1 (XNOR_1_6_N10_PULSESHAPING_OUT), .A2 (GND));

      wire XNOR_1_1_N13_PULSESHAPING_OUT, XNOR_1_2_N13_PULSESHAPING_OUT, XNOR_1_3_N13_PULSESHAPING_OUT, XNOR_1_4_N13_PULSESHAPING_OUT, XNOR_1_5_N13_PULSESHAPING_OUT, XNOR_1_6_N13_PULSESHAPING_OUT;
      NOR2_X1 XNOR_1_1_N13_PULSESHAPING (.ZN (XNOR_1_1_N13_PULSESHAPING_OUT), .A1 (N13_PWL), .A2 (GND));
      NOR2_X1 XNOR_1_2_N13_PULSESHAPING (.ZN (XNOR_1_2_N13_PULSESHAPING_OUT), .A1 (XNOR_1_1_N13_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_3_N13_PULSESHAPING (.ZN (XNOR_1_3_N13_PULSESHAPING_OUT), .A1 (XNOR_1_2_N13_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_4_N13_PULSESHAPING (.ZN (XNOR_1_4_N13_PULSESHAPING_OUT), .A1 (XNOR_1_3_N13_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_5_N13_PULSESHAPING (.ZN (XNOR_1_5_N13_PULSESHAPING_OUT), .A1 (XNOR_1_4_N13_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_6_N13_PULSESHAPING (.ZN (XNOR_1_6_N13_PULSESHAPING_OUT), .A1 (XNOR_1_5_N13_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_7_N13_PULSESHAPING (.ZN (N13), .A1 (XNOR_1_6_N13_PULSESHAPING_OUT), .A2 (GND));

      wire XNOR_1_1_N16_PULSESHAPING_OUT, XNOR_1_2_N16_PULSESHAPING_OUT, XNOR_1_3_N16_PULSESHAPING_OUT, XNOR_1_4_N16_PULSESHAPING_OUT, XNOR_1_5_N16_PULSESHAPING_OUT, XNOR_1_6_N16_PULSESHAPING_OUT;
      NOR2_X1 XNOR_1_1_N16_PULSESHAPING (.ZN (XNOR_1_1_N16_PULSESHAPING_OUT), .A1 (N16_PWL), .A2 (GND));
      NOR2_X1 XNOR_1_2_N16_PULSESHAPING (.ZN (XNOR_1_2_N16_PULSESHAPING_OUT), .A1 (XNOR_1_1_N16_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_3_N16_PULSESHAPING (.ZN (XNOR_1_3_N16_PULSESHAPING_OUT), .A1 (XNOR_1_2_N16_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_4_N16_PULSESHAPING (.ZN (XNOR_1_4_N16_PULSESHAPING_OUT), .A1 (XNOR_1_3_N16_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_5_N16_PULSESHAPING (.ZN (XNOR_1_5_N16_PULSESHAPING_OUT), .A1 (XNOR_1_4_N16_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_6_N16_PULSESHAPING (.ZN (XNOR_1_6_N16_PULSESHAPING_OUT), .A1 (XNOR_1_5_N16_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_7_N16_PULSESHAPING (.ZN (N16), .A1 (XNOR_1_6_N16_PULSESHAPING_OUT), .A2 (GND));

      wire XNOR_1_1_N19_PULSESHAPING_OUT, XNOR_1_2_N19_PULSESHAPING_OUT, XNOR_1_3_N19_PULSESHAPING_OUT, XNOR_1_4_N19_PULSESHAPING_OUT, XNOR_1_5_N19_PULSESHAPING_OUT, XNOR_1_6_N19_PULSESHAPING_OUT;
      NOR2_X1 XNOR_1_1_N19_PULSESHAPING (.ZN (XNOR_1_1_N19_PULSESHAPING_OUT), .A1 (N19_PWL), .A2 (GND));
      NOR2_X1 XNOR_1_2_N19_PULSESHAPING (.ZN (XNOR_1_2_N19_PULSESHAPING_OUT), .A1 (XNOR_1_1_N19_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_3_N19_PULSESHAPING (.ZN (XNOR_1_3_N19_PULSESHAPING_OUT), .A1 (XNOR_1_2_N19_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_4_N19_PULSESHAPING (.ZN (XNOR_1_4_N19_PULSESHAPING_OUT), .A1 (XNOR_1_3_N19_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_5_N19_PULSESHAPING (.ZN (XNOR_1_5_N19_PULSESHAPING_OUT), .A1 (XNOR_1_4_N19_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_6_N19_PULSESHAPING (.ZN (XNOR_1_6_N19_PULSESHAPING_OUT), .A1 (XNOR_1_5_N19_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_7_N19_PULSESHAPING (.ZN (N19), .A1 (XNOR_1_6_N19_PULSESHAPING_OUT), .A2 (GND));

      wire XNOR_1_1_N22_PULSESHAPING_OUT, XNOR_1_2_N22_PULSESHAPING_OUT, XNOR_1_3_N22_PULSESHAPING_OUT, XNOR_1_4_N22_PULSESHAPING_OUT, XNOR_1_5_N22_PULSESHAPING_OUT, XNOR_1_6_N22_PULSESHAPING_OUT;
      NOR2_X1 XNOR_1_1_N22_PULSESHAPING (.ZN (XNOR_1_1_N22_PULSESHAPING_OUT), .A1 (N22_PWL), .A2 (GND));
      NOR2_X1 XNOR_1_2_N22_PULSESHAPING (.ZN (XNOR_1_2_N22_PULSESHAPING_OUT), .A1 (XNOR_1_1_N22_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_3_N22_PULSESHAPING (.ZN (XNOR_1_3_N22_PULSESHAPING_OUT), .A1 (XNOR_1_2_N22_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_4_N22_PULSESHAPING (.ZN (XNOR_1_4_N22_PULSESHAPING_OUT), .A1 (XNOR_1_3_N22_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_5_N22_PULSESHAPING (.ZN (XNOR_1_5_N22_PULSESHAPING_OUT), .A1 (XNOR_1_4_N22_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_6_N22_PULSESHAPING (.ZN (XNOR_1_6_N22_PULSESHAPING_OUT), .A1 (XNOR_1_5_N22_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_7_N22_PULSESHAPING (.ZN (N22), .A1 (XNOR_1_6_N22_PULSESHAPING_OUT), .A2 (GND));

      wire XNOR_1_1_N25_PULSESHAPING_OUT, XNOR_1_2_N25_PULSESHAPING_OUT, XNOR_1_3_N25_PULSESHAPING_OUT, XNOR_1_4_N25_PULSESHAPING_OUT, XNOR_1_5_N25_PULSESHAPING_OUT, XNOR_1_6_N25_PULSESHAPING_OUT;
      NOR2_X1 XNOR_1_1_N25_PULSESHAPING (.ZN (XNOR_1_1_N25_PULSESHAPING_OUT), .A1 (N25_PWL), .A2 (GND));
      NOR2_X1 XNOR_1_2_N25_PULSESHAPING (.ZN (XNOR_1_2_N25_PULSESHAPING_OUT), .A1 (XNOR_1_1_N25_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_3_N25_PULSESHAPING (.ZN (XNOR_1_3_N25_PULSESHAPING_OUT), .A1 (XNOR_1_2_N25_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_4_N25_PULSESHAPING (.ZN (XNOR_1_4_N25_PULSESHAPING_OUT), .A1 (XNOR_1_3_N25_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_5_N25_PULSESHAPING (.ZN (XNOR_1_5_N25_PULSESHAPING_OUT), .A1 (XNOR_1_4_N25_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_6_N25_PULSESHAPING (.ZN (XNOR_1_6_N25_PULSESHAPING_OUT), .A1 (XNOR_1_5_N25_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_7_N25_PULSESHAPING (.ZN (N25), .A1 (XNOR_1_6_N25_PULSESHAPING_OUT), .A2 (GND));

      wire XNOR_1_1_N28_PULSESHAPING_OUT, XNOR_1_2_N28_PULSESHAPING_OUT, XNOR_1_3_N28_PULSESHAPING_OUT, XNOR_1_4_N28_PULSESHAPING_OUT, XNOR_1_5_N28_PULSESHAPING_OUT, XNOR_1_6_N28_PULSESHAPING_OUT;
      NOR2_X1 XNOR_1_1_N28_PULSESHAPING (.ZN (XNOR_1_1_N28_PULSESHAPING_OUT), .A1 (N28_PWL), .A2 (GND));
      NOR2_X1 XNOR_1_2_N28_PULSESHAPING (.ZN (XNOR_1_2_N28_PULSESHAPING_OUT), .A1 (XNOR_1_1_N28_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_3_N28_PULSESHAPING (.ZN (XNOR_1_3_N28_PULSESHAPING_OUT), .A1 (XNOR_1_2_N28_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_4_N28_PULSESHAPING (.ZN (XNOR_1_4_N28_PULSESHAPING_OUT), .A1 (XNOR_1_3_N28_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_5_N28_PULSESHAPING (.ZN (XNOR_1_5_N28_PULSESHAPING_OUT), .A1 (XNOR_1_4_N28_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_6_N28_PULSESHAPING (.ZN (XNOR_1_6_N28_PULSESHAPING_OUT), .A1 (XNOR_1_5_N28_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_7_N28_PULSESHAPING (.ZN (N28), .A1 (XNOR_1_6_N28_PULSESHAPING_OUT), .A2 (GND));

      wire XNOR_1_1_N31_PULSESHAPING_OUT, XNOR_1_2_N31_PULSESHAPING_OUT, XNOR_1_3_N31_PULSESHAPING_OUT, XNOR_1_4_N31_PULSESHAPING_OUT, XNOR_1_5_N31_PULSESHAPING_OUT, XNOR_1_6_N31_PULSESHAPING_OUT;
      NOR2_X1 XNOR_1_1_N31_PULSESHAPING (.ZN (XNOR_1_1_N31_PULSESHAPING_OUT), .A1 (N31_PWL), .A2 (GND));
      NOR2_X1 XNOR_1_2_N31_PULSESHAPING (.ZN (XNOR_1_2_N31_PULSESHAPING_OUT), .A1 (XNOR_1_1_N31_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_3_N31_PULSESHAPING (.ZN (XNOR_1_3_N31_PULSESHAPING_OUT), .A1 (XNOR_1_2_N31_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_4_N31_PULSESHAPING (.ZN (XNOR_1_4_N31_PULSESHAPING_OUT), .A1 (XNOR_1_3_N31_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_5_N31_PULSESHAPING (.ZN (XNOR_1_5_N31_PULSESHAPING_OUT), .A1 (XNOR_1_4_N31_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_6_N31_PULSESHAPING (.ZN (XNOR_1_6_N31_PULSESHAPING_OUT), .A1 (XNOR_1_5_N31_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_7_N31_PULSESHAPING (.ZN (N31), .A1 (XNOR_1_6_N31_PULSESHAPING_OUT), .A2 (GND));

      wire XNOR_1_1_N34_PULSESHAPING_OUT, XNOR_1_2_N34_PULSESHAPING_OUT, XNOR_1_3_N34_PULSESHAPING_OUT, XNOR_1_4_N34_PULSESHAPING_OUT, XNOR_1_5_N34_PULSESHAPING_OUT, XNOR_1_6_N34_PULSESHAPING_OUT;
      NOR2_X1 XNOR_1_1_N34_PULSESHAPING (.ZN (XNOR_1_1_N34_PULSESHAPING_OUT), .A1 (N34_PWL), .A2 (GND));
      NOR2_X1 XNOR_1_2_N34_PULSESHAPING (.ZN (XNOR_1_2_N34_PULSESHAPING_OUT), .A1 (XNOR_1_1_N34_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_3_N34_PULSESHAPING (.ZN (XNOR_1_3_N34_PULSESHAPING_OUT), .A1 (XNOR_1_2_N34_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_4_N34_PULSESHAPING (.ZN (XNOR_1_4_N34_PULSESHAPING_OUT), .A1 (XNOR_1_3_N34_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_5_N34_PULSESHAPING (.ZN (XNOR_1_5_N34_PULSESHAPING_OUT), .A1 (XNOR_1_4_N34_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_6_N34_PULSESHAPING (.ZN (XNOR_1_6_N34_PULSESHAPING_OUT), .A1 (XNOR_1_5_N34_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_7_N34_PULSESHAPING (.ZN (N34), .A1 (XNOR_1_6_N34_PULSESHAPING_OUT), .A2 (GND));

      wire XNOR_1_1_N37_PULSESHAPING_OUT, XNOR_1_2_N37_PULSESHAPING_OUT, XNOR_1_3_N37_PULSESHAPING_OUT, XNOR_1_4_N37_PULSESHAPING_OUT, XNOR_1_5_N37_PULSESHAPING_OUT, XNOR_1_6_N37_PULSESHAPING_OUT;
      NOR2_X1 XNOR_1_1_N37_PULSESHAPING (.ZN (XNOR_1_1_N37_PULSESHAPING_OUT), .A1 (N37_PWL), .A2 (GND));
      NOR2_X1 XNOR_1_2_N37_PULSESHAPING (.ZN (XNOR_1_2_N37_PULSESHAPING_OUT), .A1 (XNOR_1_1_N37_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_3_N37_PULSESHAPING (.ZN (XNOR_1_3_N37_PULSESHAPING_OUT), .A1 (XNOR_1_2_N37_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_4_N37_PULSESHAPING (.ZN (XNOR_1_4_N37_PULSESHAPING_OUT), .A1 (XNOR_1_3_N37_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_5_N37_PULSESHAPING (.ZN (XNOR_1_5_N37_PULSESHAPING_OUT), .A1 (XNOR_1_4_N37_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_6_N37_PULSESHAPING (.ZN (XNOR_1_6_N37_PULSESHAPING_OUT), .A1 (XNOR_1_5_N37_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_7_N37_PULSESHAPING (.ZN (N37), .A1 (XNOR_1_6_N37_PULSESHAPING_OUT), .A2 (GND));

      wire XNOR_1_1_N40_PULSESHAPING_OUT, XNOR_1_2_N40_PULSESHAPING_OUT, XNOR_1_3_N40_PULSESHAPING_OUT, XNOR_1_4_N40_PULSESHAPING_OUT, XNOR_1_5_N40_PULSESHAPING_OUT, XNOR_1_6_N40_PULSESHAPING_OUT;
      NOR2_X1 XNOR_1_1_N40_PULSESHAPING (.ZN (XNOR_1_1_N40_PULSESHAPING_OUT), .A1 (N40_PWL), .A2 (GND));
      NOR2_X1 XNOR_1_2_N40_PULSESHAPING (.ZN (XNOR_1_2_N40_PULSESHAPING_OUT), .A1 (XNOR_1_1_N40_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_3_N40_PULSESHAPING (.ZN (XNOR_1_3_N40_PULSESHAPING_OUT), .A1 (XNOR_1_2_N40_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_4_N40_PULSESHAPING (.ZN (XNOR_1_4_N40_PULSESHAPING_OUT), .A1 (XNOR_1_3_N40_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_5_N40_PULSESHAPING (.ZN (XNOR_1_5_N40_PULSESHAPING_OUT), .A1 (XNOR_1_4_N40_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_6_N40_PULSESHAPING (.ZN (XNOR_1_6_N40_PULSESHAPING_OUT), .A1 (XNOR_1_5_N40_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_7_N40_PULSESHAPING (.ZN (N40), .A1 (XNOR_1_6_N40_PULSESHAPING_OUT), .A2 (GND));

      wire XNOR_1_1_N43_PULSESHAPING_OUT, XNOR_1_2_N43_PULSESHAPING_OUT, XNOR_1_3_N43_PULSESHAPING_OUT, XNOR_1_4_N43_PULSESHAPING_OUT, XNOR_1_5_N43_PULSESHAPING_OUT, XNOR_1_6_N43_PULSESHAPING_OUT;
      NOR2_X1 XNOR_1_1_N43_PULSESHAPING (.ZN (XNOR_1_1_N43_PULSESHAPING_OUT), .A1 (N43_PWL), .A2 (GND));
      NOR2_X1 XNOR_1_2_N43_PULSESHAPING (.ZN (XNOR_1_2_N43_PULSESHAPING_OUT), .A1 (XNOR_1_1_N43_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_3_N43_PULSESHAPING (.ZN (XNOR_1_3_N43_PULSESHAPING_OUT), .A1 (XNOR_1_2_N43_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_4_N43_PULSESHAPING (.ZN (XNOR_1_4_N43_PULSESHAPING_OUT), .A1 (XNOR_1_3_N43_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_5_N43_PULSESHAPING (.ZN (XNOR_1_5_N43_PULSESHAPING_OUT), .A1 (XNOR_1_4_N43_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_6_N43_PULSESHAPING (.ZN (XNOR_1_6_N43_PULSESHAPING_OUT), .A1 (XNOR_1_5_N43_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_7_N43_PULSESHAPING (.ZN (N43), .A1 (XNOR_1_6_N43_PULSESHAPING_OUT), .A2 (GND));

      wire XNOR_1_1_N46_PULSESHAPING_OUT, XNOR_1_2_N46_PULSESHAPING_OUT, XNOR_1_3_N46_PULSESHAPING_OUT, XNOR_1_4_N46_PULSESHAPING_OUT, XNOR_1_5_N46_PULSESHAPING_OUT, XNOR_1_6_N46_PULSESHAPING_OUT;
      NOR2_X1 XNOR_1_1_N46_PULSESHAPING (.ZN (XNOR_1_1_N46_PULSESHAPING_OUT), .A1 (N46_PWL), .A2 (GND));
      NOR2_X1 XNOR_1_2_N46_PULSESHAPING (.ZN (XNOR_1_2_N46_PULSESHAPING_OUT), .A1 (XNOR_1_1_N46_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_3_N46_PULSESHAPING (.ZN (XNOR_1_3_N46_PULSESHAPING_OUT), .A1 (XNOR_1_2_N46_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_4_N46_PULSESHAPING (.ZN (XNOR_1_4_N46_PULSESHAPING_OUT), .A1 (XNOR_1_3_N46_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_5_N46_PULSESHAPING (.ZN (XNOR_1_5_N46_PULSESHAPING_OUT), .A1 (XNOR_1_4_N46_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_6_N46_PULSESHAPING (.ZN (XNOR_1_6_N46_PULSESHAPING_OUT), .A1 (XNOR_1_5_N46_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_7_N46_PULSESHAPING (.ZN (N46), .A1 (XNOR_1_6_N46_PULSESHAPING_OUT), .A2 (GND));

      wire XNOR_1_1_N49_PULSESHAPING_OUT, XNOR_1_2_N49_PULSESHAPING_OUT, XNOR_1_3_N49_PULSESHAPING_OUT, XNOR_1_4_N49_PULSESHAPING_OUT, XNOR_1_5_N49_PULSESHAPING_OUT, XNOR_1_6_N49_PULSESHAPING_OUT;
      NOR2_X1 XNOR_1_1_N49_PULSESHAPING (.ZN (XNOR_1_1_N49_PULSESHAPING_OUT), .A1 (N49_PWL), .A2 (GND));
      NOR2_X1 XNOR_1_2_N49_PULSESHAPING (.ZN (XNOR_1_2_N49_PULSESHAPING_OUT), .A1 (XNOR_1_1_N49_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_3_N49_PULSESHAPING (.ZN (XNOR_1_3_N49_PULSESHAPING_OUT), .A1 (XNOR_1_2_N49_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_4_N49_PULSESHAPING (.ZN (XNOR_1_4_N49_PULSESHAPING_OUT), .A1 (XNOR_1_3_N49_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_5_N49_PULSESHAPING (.ZN (XNOR_1_5_N49_PULSESHAPING_OUT), .A1 (XNOR_1_4_N49_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_6_N49_PULSESHAPING (.ZN (XNOR_1_6_N49_PULSESHAPING_OUT), .A1 (XNOR_1_5_N49_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_7_N49_PULSESHAPING (.ZN (N49), .A1 (XNOR_1_6_N49_PULSESHAPING_OUT), .A2 (GND));

      wire XNOR_1_1_N53_PULSESHAPING_OUT, XNOR_1_2_N53_PULSESHAPING_OUT, XNOR_1_3_N53_PULSESHAPING_OUT, XNOR_1_4_N53_PULSESHAPING_OUT, XNOR_1_5_N53_PULSESHAPING_OUT, XNOR_1_6_N53_PULSESHAPING_OUT;
      NOR2_X1 XNOR_1_1_N53_PULSESHAPING (.ZN (XNOR_1_1_N53_PULSESHAPING_OUT), .A1 (N53_PWL), .A2 (GND));
      NOR2_X1 XNOR_1_2_N53_PULSESHAPING (.ZN (XNOR_1_2_N53_PULSESHAPING_OUT), .A1 (XNOR_1_1_N53_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_3_N53_PULSESHAPING (.ZN (XNOR_1_3_N53_PULSESHAPING_OUT), .A1 (XNOR_1_2_N53_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_4_N53_PULSESHAPING (.ZN (XNOR_1_4_N53_PULSESHAPING_OUT), .A1 (XNOR_1_3_N53_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_5_N53_PULSESHAPING (.ZN (XNOR_1_5_N53_PULSESHAPING_OUT), .A1 (XNOR_1_4_N53_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_6_N53_PULSESHAPING (.ZN (XNOR_1_6_N53_PULSESHAPING_OUT), .A1 (XNOR_1_5_N53_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_7_N53_PULSESHAPING (.ZN (N53), .A1 (XNOR_1_6_N53_PULSESHAPING_OUT), .A2 (GND));

      wire XNOR_1_1_N56_PULSESHAPING_OUT, XNOR_1_2_N56_PULSESHAPING_OUT, XNOR_1_3_N56_PULSESHAPING_OUT, XNOR_1_4_N56_PULSESHAPING_OUT, XNOR_1_5_N56_PULSESHAPING_OUT, XNOR_1_6_N56_PULSESHAPING_OUT;
      NOR2_X1 XNOR_1_1_N56_PULSESHAPING (.ZN (XNOR_1_1_N56_PULSESHAPING_OUT), .A1 (N56_PWL), .A2 (GND));
      NOR2_X1 XNOR_1_2_N56_PULSESHAPING (.ZN (XNOR_1_2_N56_PULSESHAPING_OUT), .A1 (XNOR_1_1_N56_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_3_N56_PULSESHAPING (.ZN (XNOR_1_3_N56_PULSESHAPING_OUT), .A1 (XNOR_1_2_N56_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_4_N56_PULSESHAPING (.ZN (XNOR_1_4_N56_PULSESHAPING_OUT), .A1 (XNOR_1_3_N56_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_5_N56_PULSESHAPING (.ZN (XNOR_1_5_N56_PULSESHAPING_OUT), .A1 (XNOR_1_4_N56_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_6_N56_PULSESHAPING (.ZN (XNOR_1_6_N56_PULSESHAPING_OUT), .A1 (XNOR_1_5_N56_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_7_N56_PULSESHAPING (.ZN (N56), .A1 (XNOR_1_6_N56_PULSESHAPING_OUT), .A2 (GND));

      wire XNOR_1_1_N60_PULSESHAPING_OUT, XNOR_1_2_N60_PULSESHAPING_OUT, XNOR_1_3_N60_PULSESHAPING_OUT, XNOR_1_4_N60_PULSESHAPING_OUT, XNOR_1_5_N60_PULSESHAPING_OUT, XNOR_1_6_N60_PULSESHAPING_OUT;
      NOR2_X1 XNOR_1_1_N60_PULSESHAPING (.ZN (XNOR_1_1_N60_PULSESHAPING_OUT), .A1 (N60_PWL), .A2 (GND));
      NOR2_X1 XNOR_1_2_N60_PULSESHAPING (.ZN (XNOR_1_2_N60_PULSESHAPING_OUT), .A1 (XNOR_1_1_N60_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_3_N60_PULSESHAPING (.ZN (XNOR_1_3_N60_PULSESHAPING_OUT), .A1 (XNOR_1_2_N60_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_4_N60_PULSESHAPING (.ZN (XNOR_1_4_N60_PULSESHAPING_OUT), .A1 (XNOR_1_3_N60_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_5_N60_PULSESHAPING (.ZN (XNOR_1_5_N60_PULSESHAPING_OUT), .A1 (XNOR_1_4_N60_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_6_N60_PULSESHAPING (.ZN (XNOR_1_6_N60_PULSESHAPING_OUT), .A1 (XNOR_1_5_N60_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_7_N60_PULSESHAPING (.ZN (N60), .A1 (XNOR_1_6_N60_PULSESHAPING_OUT), .A2 (GND));

      wire XNOR_1_1_N63_PULSESHAPING_OUT, XNOR_1_2_N63_PULSESHAPING_OUT, XNOR_1_3_N63_PULSESHAPING_OUT, XNOR_1_4_N63_PULSESHAPING_OUT, XNOR_1_5_N63_PULSESHAPING_OUT, XNOR_1_6_N63_PULSESHAPING_OUT;
      NOR2_X1 XNOR_1_1_N63_PULSESHAPING (.ZN (XNOR_1_1_N63_PULSESHAPING_OUT), .A1 (N63_PWL), .A2 (GND));
      NOR2_X1 XNOR_1_2_N63_PULSESHAPING (.ZN (XNOR_1_2_N63_PULSESHAPING_OUT), .A1 (XNOR_1_1_N63_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_3_N63_PULSESHAPING (.ZN (XNOR_1_3_N63_PULSESHAPING_OUT), .A1 (XNOR_1_2_N63_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_4_N63_PULSESHAPING (.ZN (XNOR_1_4_N63_PULSESHAPING_OUT), .A1 (XNOR_1_3_N63_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_5_N63_PULSESHAPING (.ZN (XNOR_1_5_N63_PULSESHAPING_OUT), .A1 (XNOR_1_4_N63_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_6_N63_PULSESHAPING (.ZN (XNOR_1_6_N63_PULSESHAPING_OUT), .A1 (XNOR_1_5_N63_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_7_N63_PULSESHAPING (.ZN (N63), .A1 (XNOR_1_6_N63_PULSESHAPING_OUT), .A2 (GND));

      wire XNOR_1_1_N66_PULSESHAPING_OUT, XNOR_1_2_N66_PULSESHAPING_OUT, XNOR_1_3_N66_PULSESHAPING_OUT, XNOR_1_4_N66_PULSESHAPING_OUT, XNOR_1_5_N66_PULSESHAPING_OUT, XNOR_1_6_N66_PULSESHAPING_OUT;
      NOR2_X1 XNOR_1_1_N66_PULSESHAPING (.ZN (XNOR_1_1_N66_PULSESHAPING_OUT), .A1 (N66_PWL), .A2 (GND));
      NOR2_X1 XNOR_1_2_N66_PULSESHAPING (.ZN (XNOR_1_2_N66_PULSESHAPING_OUT), .A1 (XNOR_1_1_N66_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_3_N66_PULSESHAPING (.ZN (XNOR_1_3_N66_PULSESHAPING_OUT), .A1 (XNOR_1_2_N66_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_4_N66_PULSESHAPING (.ZN (XNOR_1_4_N66_PULSESHAPING_OUT), .A1 (XNOR_1_3_N66_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_5_N66_PULSESHAPING (.ZN (XNOR_1_5_N66_PULSESHAPING_OUT), .A1 (XNOR_1_4_N66_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_6_N66_PULSESHAPING (.ZN (XNOR_1_6_N66_PULSESHAPING_OUT), .A1 (XNOR_1_5_N66_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_7_N66_PULSESHAPING (.ZN (N66), .A1 (XNOR_1_6_N66_PULSESHAPING_OUT), .A2 (GND));

      wire XNOR_1_1_N69_PULSESHAPING_OUT, XNOR_1_2_N69_PULSESHAPING_OUT, XNOR_1_3_N69_PULSESHAPING_OUT, XNOR_1_4_N69_PULSESHAPING_OUT, XNOR_1_5_N69_PULSESHAPING_OUT, XNOR_1_6_N69_PULSESHAPING_OUT;
      NOR2_X1 XNOR_1_1_N69_PULSESHAPING (.ZN (XNOR_1_1_N69_PULSESHAPING_OUT), .A1 (N69_PWL), .A2 (GND));
      NOR2_X1 XNOR_1_2_N69_PULSESHAPING (.ZN (XNOR_1_2_N69_PULSESHAPING_OUT), .A1 (XNOR_1_1_N69_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_3_N69_PULSESHAPING (.ZN (XNOR_1_3_N69_PULSESHAPING_OUT), .A1 (XNOR_1_2_N69_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_4_N69_PULSESHAPING (.ZN (XNOR_1_4_N69_PULSESHAPING_OUT), .A1 (XNOR_1_3_N69_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_5_N69_PULSESHAPING (.ZN (XNOR_1_5_N69_PULSESHAPING_OUT), .A1 (XNOR_1_4_N69_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_6_N69_PULSESHAPING (.ZN (XNOR_1_6_N69_PULSESHAPING_OUT), .A1 (XNOR_1_5_N69_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_7_N69_PULSESHAPING (.ZN (N69), .A1 (XNOR_1_6_N69_PULSESHAPING_OUT), .A2 (GND));

      wire XNOR_1_1_N72_PULSESHAPING_OUT, XNOR_1_2_N72_PULSESHAPING_OUT, XNOR_1_3_N72_PULSESHAPING_OUT, XNOR_1_4_N72_PULSESHAPING_OUT, XNOR_1_5_N72_PULSESHAPING_OUT, XNOR_1_6_N72_PULSESHAPING_OUT;
      NOR2_X1 XNOR_1_1_N72_PULSESHAPING (.ZN (XNOR_1_1_N72_PULSESHAPING_OUT), .A1 (N72_PWL), .A2 (GND));
      NOR2_X1 XNOR_1_2_N72_PULSESHAPING (.ZN (XNOR_1_2_N72_PULSESHAPING_OUT), .A1 (XNOR_1_1_N72_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_3_N72_PULSESHAPING (.ZN (XNOR_1_3_N72_PULSESHAPING_OUT), .A1 (XNOR_1_2_N72_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_4_N72_PULSESHAPING (.ZN (XNOR_1_4_N72_PULSESHAPING_OUT), .A1 (XNOR_1_3_N72_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_5_N72_PULSESHAPING (.ZN (XNOR_1_5_N72_PULSESHAPING_OUT), .A1 (XNOR_1_4_N72_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_6_N72_PULSESHAPING (.ZN (XNOR_1_6_N72_PULSESHAPING_OUT), .A1 (XNOR_1_5_N72_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_7_N72_PULSESHAPING (.ZN (N72), .A1 (XNOR_1_6_N72_PULSESHAPING_OUT), .A2 (GND));

      wire XNOR_1_1_N76_PULSESHAPING_OUT, XNOR_1_2_N76_PULSESHAPING_OUT, XNOR_1_3_N76_PULSESHAPING_OUT, XNOR_1_4_N76_PULSESHAPING_OUT, XNOR_1_5_N76_PULSESHAPING_OUT, XNOR_1_6_N76_PULSESHAPING_OUT;
      NOR2_X1 XNOR_1_1_N76_PULSESHAPING (.ZN (XNOR_1_1_N76_PULSESHAPING_OUT), .A1 (N76_PWL), .A2 (GND));
      NOR2_X1 XNOR_1_2_N76_PULSESHAPING (.ZN (XNOR_1_2_N76_PULSESHAPING_OUT), .A1 (XNOR_1_1_N76_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_3_N76_PULSESHAPING (.ZN (XNOR_1_3_N76_PULSESHAPING_OUT), .A1 (XNOR_1_2_N76_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_4_N76_PULSESHAPING (.ZN (XNOR_1_4_N76_PULSESHAPING_OUT), .A1 (XNOR_1_3_N76_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_5_N76_PULSESHAPING (.ZN (XNOR_1_5_N76_PULSESHAPING_OUT), .A1 (XNOR_1_4_N76_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_6_N76_PULSESHAPING (.ZN (XNOR_1_6_N76_PULSESHAPING_OUT), .A1 (XNOR_1_5_N76_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_7_N76_PULSESHAPING (.ZN (N76), .A1 (XNOR_1_6_N76_PULSESHAPING_OUT), .A2 (GND));

      wire XNOR_1_1_N79_PULSESHAPING_OUT, XNOR_1_2_N79_PULSESHAPING_OUT, XNOR_1_3_N79_PULSESHAPING_OUT, XNOR_1_4_N79_PULSESHAPING_OUT, XNOR_1_5_N79_PULSESHAPING_OUT, XNOR_1_6_N79_PULSESHAPING_OUT;
      NOR2_X1 XNOR_1_1_N79_PULSESHAPING (.ZN (XNOR_1_1_N79_PULSESHAPING_OUT), .A1 (N79_PWL), .A2 (GND));
      NOR2_X1 XNOR_1_2_N79_PULSESHAPING (.ZN (XNOR_1_2_N79_PULSESHAPING_OUT), .A1 (XNOR_1_1_N79_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_3_N79_PULSESHAPING (.ZN (XNOR_1_3_N79_PULSESHAPING_OUT), .A1 (XNOR_1_2_N79_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_4_N79_PULSESHAPING (.ZN (XNOR_1_4_N79_PULSESHAPING_OUT), .A1 (XNOR_1_3_N79_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_5_N79_PULSESHAPING (.ZN (XNOR_1_5_N79_PULSESHAPING_OUT), .A1 (XNOR_1_4_N79_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_6_N79_PULSESHAPING (.ZN (XNOR_1_6_N79_PULSESHAPING_OUT), .A1 (XNOR_1_5_N79_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_7_N79_PULSESHAPING (.ZN (N79), .A1 (XNOR_1_6_N79_PULSESHAPING_OUT), .A2 (GND));

      wire XNOR_1_1_N82_PULSESHAPING_OUT, XNOR_1_2_N82_PULSESHAPING_OUT, XNOR_1_3_N82_PULSESHAPING_OUT, XNOR_1_4_N82_PULSESHAPING_OUT, XNOR_1_5_N82_PULSESHAPING_OUT, XNOR_1_6_N82_PULSESHAPING_OUT;
      NOR2_X1 XNOR_1_1_N82_PULSESHAPING (.ZN (XNOR_1_1_N82_PULSESHAPING_OUT), .A1 (N82_PWL), .A2 (GND));
      NOR2_X1 XNOR_1_2_N82_PULSESHAPING (.ZN (XNOR_1_2_N82_PULSESHAPING_OUT), .A1 (XNOR_1_1_N82_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_3_N82_PULSESHAPING (.ZN (XNOR_1_3_N82_PULSESHAPING_OUT), .A1 (XNOR_1_2_N82_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_4_N82_PULSESHAPING (.ZN (XNOR_1_4_N82_PULSESHAPING_OUT), .A1 (XNOR_1_3_N82_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_5_N82_PULSESHAPING (.ZN (XNOR_1_5_N82_PULSESHAPING_OUT), .A1 (XNOR_1_4_N82_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_6_N82_PULSESHAPING (.ZN (XNOR_1_6_N82_PULSESHAPING_OUT), .A1 (XNOR_1_5_N82_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_7_N82_PULSESHAPING (.ZN (N82), .A1 (XNOR_1_6_N82_PULSESHAPING_OUT), .A2 (GND));

      wire XNOR_1_1_N85_PULSESHAPING_OUT, XNOR_1_2_N85_PULSESHAPING_OUT, XNOR_1_3_N85_PULSESHAPING_OUT, XNOR_1_4_N85_PULSESHAPING_OUT, XNOR_1_5_N85_PULSESHAPING_OUT, XNOR_1_6_N85_PULSESHAPING_OUT;
      NOR2_X1 XNOR_1_1_N85_PULSESHAPING (.ZN (XNOR_1_1_N85_PULSESHAPING_OUT), .A1 (N85_PWL), .A2 (GND));
      NOR2_X1 XNOR_1_2_N85_PULSESHAPING (.ZN (XNOR_1_2_N85_PULSESHAPING_OUT), .A1 (XNOR_1_1_N85_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_3_N85_PULSESHAPING (.ZN (XNOR_1_3_N85_PULSESHAPING_OUT), .A1 (XNOR_1_2_N85_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_4_N85_PULSESHAPING (.ZN (XNOR_1_4_N85_PULSESHAPING_OUT), .A1 (XNOR_1_3_N85_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_5_N85_PULSESHAPING (.ZN (XNOR_1_5_N85_PULSESHAPING_OUT), .A1 (XNOR_1_4_N85_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_6_N85_PULSESHAPING (.ZN (XNOR_1_6_N85_PULSESHAPING_OUT), .A1 (XNOR_1_5_N85_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_7_N85_PULSESHAPING (.ZN (N85), .A1 (XNOR_1_6_N85_PULSESHAPING_OUT), .A2 (GND));

      wire XNOR_1_1_N88_PULSESHAPING_OUT, XNOR_1_2_N88_PULSESHAPING_OUT, XNOR_1_3_N88_PULSESHAPING_OUT, XNOR_1_4_N88_PULSESHAPING_OUT, XNOR_1_5_N88_PULSESHAPING_OUT, XNOR_1_6_N88_PULSESHAPING_OUT;
      NOR2_X1 XNOR_1_1_N88_PULSESHAPING (.ZN (XNOR_1_1_N88_PULSESHAPING_OUT), .A1 (N88_PWL), .A2 (GND));
      NOR2_X1 XNOR_1_2_N88_PULSESHAPING (.ZN (XNOR_1_2_N88_PULSESHAPING_OUT), .A1 (XNOR_1_1_N88_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_3_N88_PULSESHAPING (.ZN (XNOR_1_3_N88_PULSESHAPING_OUT), .A1 (XNOR_1_2_N88_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_4_N88_PULSESHAPING (.ZN (XNOR_1_4_N88_PULSESHAPING_OUT), .A1 (XNOR_1_3_N88_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_5_N88_PULSESHAPING (.ZN (XNOR_1_5_N88_PULSESHAPING_OUT), .A1 (XNOR_1_4_N88_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_6_N88_PULSESHAPING (.ZN (XNOR_1_6_N88_PULSESHAPING_OUT), .A1 (XNOR_1_5_N88_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_7_N88_PULSESHAPING (.ZN (N88), .A1 (XNOR_1_6_N88_PULSESHAPING_OUT), .A2 (GND));

      wire XNOR_1_1_N91_PULSESHAPING_OUT, XNOR_1_2_N91_PULSESHAPING_OUT, XNOR_1_3_N91_PULSESHAPING_OUT, XNOR_1_4_N91_PULSESHAPING_OUT, XNOR_1_5_N91_PULSESHAPING_OUT, XNOR_1_6_N91_PULSESHAPING_OUT;
      NOR2_X1 XNOR_1_1_N91_PULSESHAPING (.ZN (XNOR_1_1_N91_PULSESHAPING_OUT), .A1 (N91_PWL), .A2 (GND));
      NOR2_X1 XNOR_1_2_N91_PULSESHAPING (.ZN (XNOR_1_2_N91_PULSESHAPING_OUT), .A1 (XNOR_1_1_N91_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_3_N91_PULSESHAPING (.ZN (XNOR_1_3_N91_PULSESHAPING_OUT), .A1 (XNOR_1_2_N91_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_4_N91_PULSESHAPING (.ZN (XNOR_1_4_N91_PULSESHAPING_OUT), .A1 (XNOR_1_3_N91_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_5_N91_PULSESHAPING (.ZN (XNOR_1_5_N91_PULSESHAPING_OUT), .A1 (XNOR_1_4_N91_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_6_N91_PULSESHAPING (.ZN (XNOR_1_6_N91_PULSESHAPING_OUT), .A1 (XNOR_1_5_N91_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_7_N91_PULSESHAPING (.ZN (N91), .A1 (XNOR_1_6_N91_PULSESHAPING_OUT), .A2 (GND));

      wire XNOR_1_1_N94_PULSESHAPING_OUT, XNOR_1_2_N94_PULSESHAPING_OUT, XNOR_1_3_N94_PULSESHAPING_OUT, XNOR_1_4_N94_PULSESHAPING_OUT, XNOR_1_5_N94_PULSESHAPING_OUT, XNOR_1_6_N94_PULSESHAPING_OUT;
      NOR2_X1 XNOR_1_1_N94_PULSESHAPING (.ZN (XNOR_1_1_N94_PULSESHAPING_OUT), .A1 (N94_PWL), .A2 (GND));
      NOR2_X1 XNOR_1_2_N94_PULSESHAPING (.ZN (XNOR_1_2_N94_PULSESHAPING_OUT), .A1 (XNOR_1_1_N94_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_3_N94_PULSESHAPING (.ZN (XNOR_1_3_N94_PULSESHAPING_OUT), .A1 (XNOR_1_2_N94_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_4_N94_PULSESHAPING (.ZN (XNOR_1_4_N94_PULSESHAPING_OUT), .A1 (XNOR_1_3_N94_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_5_N94_PULSESHAPING (.ZN (XNOR_1_5_N94_PULSESHAPING_OUT), .A1 (XNOR_1_4_N94_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_6_N94_PULSESHAPING (.ZN (XNOR_1_6_N94_PULSESHAPING_OUT), .A1 (XNOR_1_5_N94_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_7_N94_PULSESHAPING (.ZN (N94), .A1 (XNOR_1_6_N94_PULSESHAPING_OUT), .A2 (GND));

      wire XNOR_1_1_N99_PULSESHAPING_OUT, XNOR_1_2_N99_PULSESHAPING_OUT, XNOR_1_3_N99_PULSESHAPING_OUT, XNOR_1_4_N99_PULSESHAPING_OUT, XNOR_1_5_N99_PULSESHAPING_OUT, XNOR_1_6_N99_PULSESHAPING_OUT;
      NOR2_X1 XNOR_1_1_N99_PULSESHAPING (.ZN (XNOR_1_1_N99_PULSESHAPING_OUT), .A1 (N99_PWL), .A2 (GND));
      NOR2_X1 XNOR_1_2_N99_PULSESHAPING (.ZN (XNOR_1_2_N99_PULSESHAPING_OUT), .A1 (XNOR_1_1_N99_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_3_N99_PULSESHAPING (.ZN (XNOR_1_3_N99_PULSESHAPING_OUT), .A1 (XNOR_1_2_N99_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_4_N99_PULSESHAPING (.ZN (XNOR_1_4_N99_PULSESHAPING_OUT), .A1 (XNOR_1_3_N99_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_5_N99_PULSESHAPING (.ZN (XNOR_1_5_N99_PULSESHAPING_OUT), .A1 (XNOR_1_4_N99_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_6_N99_PULSESHAPING (.ZN (XNOR_1_6_N99_PULSESHAPING_OUT), .A1 (XNOR_1_5_N99_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_7_N99_PULSESHAPING (.ZN (N99), .A1 (XNOR_1_6_N99_PULSESHAPING_OUT), .A2 (GND));

      wire XNOR_1_1_N104_PULSESHAPING_OUT, XNOR_1_2_N104_PULSESHAPING_OUT, XNOR_1_3_N104_PULSESHAPING_OUT, XNOR_1_4_N104_PULSESHAPING_OUT, XNOR_1_5_N104_PULSESHAPING_OUT, XNOR_1_6_N104_PULSESHAPING_OUT;
      NOR2_X1 XNOR_1_1_N104_PULSESHAPING (.ZN (XNOR_1_1_N104_PULSESHAPING_OUT), .A1 (N104_PWL), .A2 (GND));
      NOR2_X1 XNOR_1_2_N104_PULSESHAPING (.ZN (XNOR_1_2_N104_PULSESHAPING_OUT), .A1 (XNOR_1_1_N104_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_3_N104_PULSESHAPING (.ZN (XNOR_1_3_N104_PULSESHAPING_OUT), .A1 (XNOR_1_2_N104_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_4_N104_PULSESHAPING (.ZN (XNOR_1_4_N104_PULSESHAPING_OUT), .A1 (XNOR_1_3_N104_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_5_N104_PULSESHAPING (.ZN (XNOR_1_5_N104_PULSESHAPING_OUT), .A1 (XNOR_1_4_N104_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_6_N104_PULSESHAPING (.ZN (XNOR_1_6_N104_PULSESHAPING_OUT), .A1 (XNOR_1_5_N104_PULSESHAPING_OUT), .A2 (GND));
      NOR2_X1 XNOR_1_7_N104_PULSESHAPING (.ZN (N104), .A1 (XNOR_1_6_N104_PULSESHAPING_OUT), .A2 (GND));



      NOR2_X1 XNOR_NOT1_NUM1 (.ZN (N190), .A1 (N1), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM2 (.ZN (N194), .A1 (N4), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM3 (.ZN (N197), .A1 (N7), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM4 (.ZN (N201), .A1 (N10), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM5 (.ZN (N206), .A1 (N13), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM6 (.ZN (N209), .A1 (N16), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM7 (.ZN (N212), .A1 (N19), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM8 (.ZN (N216), .A1 (N22), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM9 (.ZN (N220), .A1 (N25), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM10 (.ZN (N225), .A1 (N28), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM11 (.ZN (N229), .A1 (N31), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM12 (.ZN (N232), .A1 (N34), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM13 (.ZN (N235), .A1 (N37), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM14 (.ZN (N239), .A1 (N40), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM15 (.ZN (N243), .A1 (N43), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM16 (.ZN (N247), .A1 (N46), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM17_OUT, XNOR_1_2_NAND2_NUM17_OUT, XNOR_1_3_NAND2_NUM17_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM17 (.ZN (XNOR_1_1_NAND2_NUM17_OUT), .A1 (N63), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM17 (.ZN (XNOR_1_2_NAND2_NUM17_OUT), .A1 (GND), .A2 (N88));
      NOR2_X1 XNOR_1_3_NAND2_NUM17 (.ZN (XNOR_1_3_NAND2_NUM17_OUT), .A1 (XNOR_1_1_NAND2_NUM17_OUT), .A2 (XNOR_1_2_NAND2_NUM17_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM17 (.ZN (N251), .A1 (XNOR_1_3_NAND2_NUM17_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM18_OUT, XNOR_1_2_NAND2_NUM18_OUT, XNOR_1_3_NAND2_NUM18_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM18 (.ZN (XNOR_1_1_NAND2_NUM18_OUT), .A1 (N66), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM18 (.ZN (XNOR_1_2_NAND2_NUM18_OUT), .A1 (GND), .A2 (N91));
      NOR2_X1 XNOR_1_3_NAND2_NUM18 (.ZN (XNOR_1_3_NAND2_NUM18_OUT), .A1 (XNOR_1_1_NAND2_NUM18_OUT), .A2 (XNOR_1_2_NAND2_NUM18_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM18 (.ZN (N252), .A1 (XNOR_1_3_NAND2_NUM18_OUT), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM19 (.ZN (N253), .A1 (N72), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM20 (.ZN (N256), .A1 (N72), .A2 (GND));
      wire XNOR_1_1_BUFF1_NUM21_OUT;
      NOR2_X1 XNOR_1_1_BUFF1_NUM21 (.ZN (XNOR_1_1_BUFF1_NUM21_OUT), .A1 (N69), .A2 (GND));
      NOR2_X1 XNOR_1_2_BUFF1_NUM21 (.ZN (N257), .A1 (XNOR_1_1_BUFF1_NUM21_OUT), .A2 (GND));
      wire XNOR_1_1_BUFF1_NUM22_OUT;
      NOR2_X1 XNOR_1_1_BUFF1_NUM22 (.ZN (XNOR_1_1_BUFF1_NUM22_OUT), .A1 (N69), .A2 (GND));
      NOR2_X1 XNOR_1_2_BUFF1_NUM22 (.ZN (N260), .A1 (XNOR_1_1_BUFF1_NUM22_OUT), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM23 (.ZN (N263), .A1 (N76), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM24 (.ZN (N266), .A1 (N79), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM25 (.ZN (N269), .A1 (N82), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM26 (.ZN (N272), .A1 (N85), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM27 (.ZN (N275), .A1 (N104), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM28 (.ZN (N276), .A1 (N104), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM29 (.ZN (N277), .A1 (N88), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM30 (.ZN (N280), .A1 (N91), .A2 (GND));
      wire XNOR_1_1_BUFF1_NUM31_OUT;
      NOR2_X1 XNOR_1_1_BUFF1_NUM31 (.ZN (XNOR_1_1_BUFF1_NUM31_OUT), .A1 (N94), .A2 (GND));
      NOR2_X1 XNOR_1_2_BUFF1_NUM31 (.ZN (N283), .A1 (XNOR_1_1_BUFF1_NUM31_OUT), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM32 (.ZN (N290), .A1 (N94), .A2 (GND));
      wire XNOR_1_1_BUFF1_NUM33_OUT;
      NOR2_X1 XNOR_1_1_BUFF1_NUM33 (.ZN (XNOR_1_1_BUFF1_NUM33_OUT), .A1 (N94), .A2 (GND));
      NOR2_X1 XNOR_1_2_BUFF1_NUM33 (.ZN (N297), .A1 (XNOR_1_1_BUFF1_NUM33_OUT), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM34 (.ZN (N300), .A1 (N94), .A2 (GND));
      wire XNOR_1_1_BUFF1_NUM35_OUT;
      NOR2_X1 XNOR_1_1_BUFF1_NUM35 (.ZN (XNOR_1_1_BUFF1_NUM35_OUT), .A1 (N99), .A2 (GND));
      NOR2_X1 XNOR_1_2_BUFF1_NUM35 (.ZN (N303), .A1 (XNOR_1_1_BUFF1_NUM35_OUT), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM36 (.ZN (N306), .A1 (N99), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM37 (.ZN (N313), .A1 (N99), .A2 (GND));
      wire XNOR_1_1_BUFF1_NUM38_OUT;
      NOR2_X1 XNOR_1_1_BUFF1_NUM38 (.ZN (XNOR_1_1_BUFF1_NUM38_OUT), .A1 (N104), .A2 (GND));
      NOR2_X1 XNOR_1_2_BUFF1_NUM38 (.ZN (N316), .A1 (XNOR_1_1_BUFF1_NUM38_OUT), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM39 (.ZN (N319), .A1 (N104), .A2 (GND));
      wire XNOR_1_1_BUFF1_NUM40_OUT;
      NOR2_X1 XNOR_1_1_BUFF1_NUM40 (.ZN (XNOR_1_1_BUFF1_NUM40_OUT), .A1 (N104), .A2 (GND));
      NOR2_X1 XNOR_1_2_BUFF1_NUM40 (.ZN (N326), .A1 (XNOR_1_1_BUFF1_NUM40_OUT), .A2 (GND));
      wire XNOR_1_1_BUFF1_NUM41_OUT;
      NOR2_X1 XNOR_1_1_BUFF1_NUM41 (.ZN (XNOR_1_1_BUFF1_NUM41_OUT), .A1 (N104), .A2 (GND));
      NOR2_X1 XNOR_1_2_BUFF1_NUM41 (.ZN (N331), .A1 (XNOR_1_1_BUFF1_NUM41_OUT), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM42 (.ZN (N338), .A1 (N104), .A2 (GND));
      wire XNOR_1_1_BUFF1_NUM43_OUT;
      NOR2_X1 XNOR_1_1_BUFF1_NUM43 (.ZN (XNOR_1_1_BUFF1_NUM43_OUT), .A1 (N1), .A2 (GND));
      NOR2_X1 XNOR_1_2_BUFF1_NUM43 (.ZN (N343), .A1 (XNOR_1_1_BUFF1_NUM43_OUT), .A2 (GND));
      wire XNOR_1_1_BUFF1_NUM44_OUT;
      NOR2_X1 XNOR_1_1_BUFF1_NUM44 (.ZN (XNOR_1_1_BUFF1_NUM44_OUT), .A1 (N4), .A2 (GND));
      NOR2_X1 XNOR_1_2_BUFF1_NUM44 (.ZN (N346), .A1 (XNOR_1_1_BUFF1_NUM44_OUT), .A2 (GND));
      wire XNOR_1_1_BUFF1_NUM45_OUT;
      NOR2_X1 XNOR_1_1_BUFF1_NUM45 (.ZN (XNOR_1_1_BUFF1_NUM45_OUT), .A1 (N7), .A2 (GND));
      NOR2_X1 XNOR_1_2_BUFF1_NUM45 (.ZN (N349), .A1 (XNOR_1_1_BUFF1_NUM45_OUT), .A2 (GND));
      wire XNOR_1_1_BUFF1_NUM46_OUT;
      NOR2_X1 XNOR_1_1_BUFF1_NUM46 (.ZN (XNOR_1_1_BUFF1_NUM46_OUT), .A1 (N10), .A2 (GND));
      NOR2_X1 XNOR_1_2_BUFF1_NUM46 (.ZN (N352), .A1 (XNOR_1_1_BUFF1_NUM46_OUT), .A2 (GND));
      wire XNOR_1_1_BUFF1_NUM47_OUT;
      NOR2_X1 XNOR_1_1_BUFF1_NUM47 (.ZN (XNOR_1_1_BUFF1_NUM47_OUT), .A1 (N13), .A2 (GND));
      NOR2_X1 XNOR_1_2_BUFF1_NUM47 (.ZN (N355), .A1 (XNOR_1_1_BUFF1_NUM47_OUT), .A2 (GND));
      wire XNOR_1_1_BUFF1_NUM48_OUT;
      NOR2_X1 XNOR_1_1_BUFF1_NUM48 (.ZN (XNOR_1_1_BUFF1_NUM48_OUT), .A1 (N16), .A2 (GND));
      NOR2_X1 XNOR_1_2_BUFF1_NUM48 (.ZN (N358), .A1 (XNOR_1_1_BUFF1_NUM48_OUT), .A2 (GND));
      wire XNOR_1_1_BUFF1_NUM49_OUT;
      NOR2_X1 XNOR_1_1_BUFF1_NUM49 (.ZN (XNOR_1_1_BUFF1_NUM49_OUT), .A1 (N19), .A2 (GND));
      NOR2_X1 XNOR_1_2_BUFF1_NUM49 (.ZN (N361), .A1 (XNOR_1_1_BUFF1_NUM49_OUT), .A2 (GND));
      wire XNOR_1_1_BUFF1_NUM50_OUT;
      NOR2_X1 XNOR_1_1_BUFF1_NUM50 (.ZN (XNOR_1_1_BUFF1_NUM50_OUT), .A1 (N22), .A2 (GND));
      NOR2_X1 XNOR_1_2_BUFF1_NUM50 (.ZN (N364), .A1 (XNOR_1_1_BUFF1_NUM50_OUT), .A2 (GND));
      wire XNOR_1_1_BUFF1_NUM51_OUT;
      NOR2_X1 XNOR_1_1_BUFF1_NUM51 (.ZN (XNOR_1_1_BUFF1_NUM51_OUT), .A1 (N25), .A2 (GND));
      NOR2_X1 XNOR_1_2_BUFF1_NUM51 (.ZN (N367), .A1 (XNOR_1_1_BUFF1_NUM51_OUT), .A2 (GND));
      wire XNOR_1_1_BUFF1_NUM52_OUT;
      NOR2_X1 XNOR_1_1_BUFF1_NUM52 (.ZN (XNOR_1_1_BUFF1_NUM52_OUT), .A1 (N28), .A2 (GND));
      NOR2_X1 XNOR_1_2_BUFF1_NUM52 (.ZN (N370), .A1 (XNOR_1_1_BUFF1_NUM52_OUT), .A2 (GND));
      wire XNOR_1_1_BUFF1_NUM53_OUT;
      NOR2_X1 XNOR_1_1_BUFF1_NUM53 (.ZN (XNOR_1_1_BUFF1_NUM53_OUT), .A1 (N31), .A2 (GND));
      NOR2_X1 XNOR_1_2_BUFF1_NUM53 (.ZN (N373), .A1 (XNOR_1_1_BUFF1_NUM53_OUT), .A2 (GND));
      wire XNOR_1_1_BUFF1_NUM54_OUT;
      NOR2_X1 XNOR_1_1_BUFF1_NUM54 (.ZN (XNOR_1_1_BUFF1_NUM54_OUT), .A1 (N34), .A2 (GND));
      NOR2_X1 XNOR_1_2_BUFF1_NUM54 (.ZN (N376), .A1 (XNOR_1_1_BUFF1_NUM54_OUT), .A2 (GND));
      wire XNOR_1_1_BUFF1_NUM55_OUT;
      NOR2_X1 XNOR_1_1_BUFF1_NUM55 (.ZN (XNOR_1_1_BUFF1_NUM55_OUT), .A1 (N37), .A2 (GND));
      NOR2_X1 XNOR_1_2_BUFF1_NUM55 (.ZN (N379), .A1 (XNOR_1_1_BUFF1_NUM55_OUT), .A2 (GND));
      wire XNOR_1_1_BUFF1_NUM56_OUT;
      NOR2_X1 XNOR_1_1_BUFF1_NUM56 (.ZN (XNOR_1_1_BUFF1_NUM56_OUT), .A1 (N40), .A2 (GND));
      NOR2_X1 XNOR_1_2_BUFF1_NUM56 (.ZN (N382), .A1 (XNOR_1_1_BUFF1_NUM56_OUT), .A2 (GND));
      wire XNOR_1_1_BUFF1_NUM57_OUT;
      NOR2_X1 XNOR_1_1_BUFF1_NUM57 (.ZN (XNOR_1_1_BUFF1_NUM57_OUT), .A1 (N43), .A2 (GND));
      NOR2_X1 XNOR_1_2_BUFF1_NUM57 (.ZN (N385), .A1 (XNOR_1_1_BUFF1_NUM57_OUT), .A2 (GND));
      wire XNOR_1_1_BUFF1_NUM58_OUT;
      NOR2_X1 XNOR_1_1_BUFF1_NUM58 (.ZN (XNOR_1_1_BUFF1_NUM58_OUT), .A1 (N46), .A2 (GND));
      NOR2_X1 XNOR_1_2_BUFF1_NUM58 (.ZN (N388), .A1 (XNOR_1_1_BUFF1_NUM58_OUT), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM59 (.ZN (N534), .A1 (N343), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM60 (.ZN (N535), .A1 (N346), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM61 (.ZN (N536), .A1 (N349), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM62 (.ZN (N537), .A1 (N352), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM63 (.ZN (N538), .A1 (N355), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM64 (.ZN (N539), .A1 (N358), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM65 (.ZN (N540), .A1 (N361), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM66 (.ZN (N541), .A1 (N364), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM67 (.ZN (N542), .A1 (N367), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM68 (.ZN (N543), .A1 (N370), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM69 (.ZN (N544), .A1 (N373), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM70 (.ZN (N545), .A1 (N376), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM71 (.ZN (N546), .A1 (N379), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM72 (.ZN (N547), .A1 (N382), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM73 (.ZN (N548), .A1 (N385), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM74 (.ZN (N549), .A1 (N388), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM75_OUT, XNOR_1_2_NAND2_NUM75_OUT, XNOR_1_3_NAND2_NUM75_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM75 (.ZN (XNOR_1_1_NAND2_NUM75_OUT), .A1 (N306), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM75 (.ZN (XNOR_1_2_NAND2_NUM75_OUT), .A1 (GND), .A2 (N331));
      NOR2_X1 XNOR_1_3_NAND2_NUM75 (.ZN (XNOR_1_3_NAND2_NUM75_OUT), .A1 (XNOR_1_1_NAND2_NUM75_OUT), .A2 (XNOR_1_2_NAND2_NUM75_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM75 (.ZN (N550), .A1 (XNOR_1_3_NAND2_NUM75_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM76_OUT, XNOR_1_2_NAND2_NUM76_OUT, XNOR_1_3_NAND2_NUM76_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM76 (.ZN (XNOR_1_1_NAND2_NUM76_OUT), .A1 (N306), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM76 (.ZN (XNOR_1_2_NAND2_NUM76_OUT), .A1 (GND), .A2 (N331));
      NOR2_X1 XNOR_1_3_NAND2_NUM76 (.ZN (XNOR_1_3_NAND2_NUM76_OUT), .A1 (XNOR_1_1_NAND2_NUM76_OUT), .A2 (XNOR_1_2_NAND2_NUM76_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM76 (.ZN (N551), .A1 (XNOR_1_3_NAND2_NUM76_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM77_OUT, XNOR_1_2_NAND2_NUM77_OUT, XNOR_1_3_NAND2_NUM77_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM77 (.ZN (XNOR_1_1_NAND2_NUM77_OUT), .A1 (N306), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM77 (.ZN (XNOR_1_2_NAND2_NUM77_OUT), .A1 (GND), .A2 (N331));
      NOR2_X1 XNOR_1_3_NAND2_NUM77 (.ZN (XNOR_1_3_NAND2_NUM77_OUT), .A1 (XNOR_1_1_NAND2_NUM77_OUT), .A2 (XNOR_1_2_NAND2_NUM77_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM77 (.ZN (N552), .A1 (XNOR_1_3_NAND2_NUM77_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM78_OUT, XNOR_1_2_NAND2_NUM78_OUT, XNOR_1_3_NAND2_NUM78_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM78 (.ZN (XNOR_1_1_NAND2_NUM78_OUT), .A1 (N306), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM78 (.ZN (XNOR_1_2_NAND2_NUM78_OUT), .A1 (GND), .A2 (N331));
      NOR2_X1 XNOR_1_3_NAND2_NUM78 (.ZN (XNOR_1_3_NAND2_NUM78_OUT), .A1 (XNOR_1_1_NAND2_NUM78_OUT), .A2 (XNOR_1_2_NAND2_NUM78_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM78 (.ZN (N553), .A1 (XNOR_1_3_NAND2_NUM78_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM79_OUT, XNOR_1_2_NAND2_NUM79_OUT, XNOR_1_3_NAND2_NUM79_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM79 (.ZN (XNOR_1_1_NAND2_NUM79_OUT), .A1 (N306), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM79 (.ZN (XNOR_1_2_NAND2_NUM79_OUT), .A1 (GND), .A2 (N331));
      NOR2_X1 XNOR_1_3_NAND2_NUM79 (.ZN (XNOR_1_3_NAND2_NUM79_OUT), .A1 (XNOR_1_1_NAND2_NUM79_OUT), .A2 (XNOR_1_2_NAND2_NUM79_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM79 (.ZN (N554), .A1 (XNOR_1_3_NAND2_NUM79_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM80_OUT, XNOR_1_2_NAND2_NUM80_OUT, XNOR_1_3_NAND2_NUM80_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM80 (.ZN (XNOR_1_1_NAND2_NUM80_OUT), .A1 (N306), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM80 (.ZN (XNOR_1_2_NAND2_NUM80_OUT), .A1 (GND), .A2 (N331));
      NOR2_X1 XNOR_1_3_NAND2_NUM80 (.ZN (XNOR_1_3_NAND2_NUM80_OUT), .A1 (XNOR_1_1_NAND2_NUM80_OUT), .A2 (XNOR_1_2_NAND2_NUM80_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM80 (.ZN (N555), .A1 (XNOR_1_3_NAND2_NUM80_OUT), .A2 (GND));
      wire XNOR_1_1_BUFF1_NUM81_OUT;
      NOR2_X1 XNOR_1_1_BUFF1_NUM81 (.ZN (XNOR_1_1_BUFF1_NUM81_OUT), .A1 (N190), .A2 (GND));
      NOR2_X1 XNOR_1_2_BUFF1_NUM81 (.ZN (N556), .A1 (XNOR_1_1_BUFF1_NUM81_OUT), .A2 (GND));
      wire XNOR_1_1_BUFF1_NUM82_OUT;
      NOR2_X1 XNOR_1_1_BUFF1_NUM82 (.ZN (XNOR_1_1_BUFF1_NUM82_OUT), .A1 (N194), .A2 (GND));
      NOR2_X1 XNOR_1_2_BUFF1_NUM82 (.ZN (N559), .A1 (XNOR_1_1_BUFF1_NUM82_OUT), .A2 (GND));
      wire XNOR_1_1_BUFF1_NUM83_OUT;
      NOR2_X1 XNOR_1_1_BUFF1_NUM83 (.ZN (XNOR_1_1_BUFF1_NUM83_OUT), .A1 (N206), .A2 (GND));
      NOR2_X1 XNOR_1_2_BUFF1_NUM83 (.ZN (N562), .A1 (XNOR_1_1_BUFF1_NUM83_OUT), .A2 (GND));
      wire XNOR_1_1_BUFF1_NUM84_OUT;
      NOR2_X1 XNOR_1_1_BUFF1_NUM84 (.ZN (XNOR_1_1_BUFF1_NUM84_OUT), .A1 (N209), .A2 (GND));
      NOR2_X1 XNOR_1_2_BUFF1_NUM84 (.ZN (N565), .A1 (XNOR_1_1_BUFF1_NUM84_OUT), .A2 (GND));
      wire XNOR_1_1_BUFF1_NUM85_OUT;
      NOR2_X1 XNOR_1_1_BUFF1_NUM85 (.ZN (XNOR_1_1_BUFF1_NUM85_OUT), .A1 (N225), .A2 (GND));
      NOR2_X1 XNOR_1_2_BUFF1_NUM85 (.ZN (N568), .A1 (XNOR_1_1_BUFF1_NUM85_OUT), .A2 (GND));
      wire XNOR_1_1_BUFF1_NUM86_OUT;
      NOR2_X1 XNOR_1_1_BUFF1_NUM86 (.ZN (XNOR_1_1_BUFF1_NUM86_OUT), .A1 (N243), .A2 (GND));
      NOR2_X1 XNOR_1_2_BUFF1_NUM86 (.ZN (N571), .A1 (XNOR_1_1_BUFF1_NUM86_OUT), .A2 (GND));
      wire XNOR_1_1_AND2_NUM87_OUT, XNOR_1_2_AND2_NUM87_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM87 (.ZN (XNOR_1_1_AND2_NUM87_OUT), .A1 (N63), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM87 (.ZN (XNOR_1_2_AND2_NUM87_OUT), .A1 (GND), .A2 (N319));
      NOR2_X1 XNOR_1_3_AND2_NUM87 (.ZN (N574), .A1 (XNOR_1_1_AND2_NUM87_OUT), .A2 (XNOR_1_2_AND2_NUM87_OUT));
      wire XNOR_1_1_BUFF1_NUM88_OUT;
      NOR2_X1 XNOR_1_1_BUFF1_NUM88 (.ZN (XNOR_1_1_BUFF1_NUM88_OUT), .A1 (N220), .A2 (GND));
      NOR2_X1 XNOR_1_2_BUFF1_NUM88 (.ZN (N577), .A1 (XNOR_1_1_BUFF1_NUM88_OUT), .A2 (GND));
      wire XNOR_1_1_BUFF1_NUM89_OUT;
      NOR2_X1 XNOR_1_1_BUFF1_NUM89 (.ZN (XNOR_1_1_BUFF1_NUM89_OUT), .A1 (N229), .A2 (GND));
      NOR2_X1 XNOR_1_2_BUFF1_NUM89 (.ZN (N580), .A1 (XNOR_1_1_BUFF1_NUM89_OUT), .A2 (GND));
      wire XNOR_1_1_BUFF1_NUM90_OUT;
      NOR2_X1 XNOR_1_1_BUFF1_NUM90 (.ZN (XNOR_1_1_BUFF1_NUM90_OUT), .A1 (N232), .A2 (GND));
      NOR2_X1 XNOR_1_2_BUFF1_NUM90 (.ZN (N583), .A1 (XNOR_1_1_BUFF1_NUM90_OUT), .A2 (GND));
      wire XNOR_1_1_AND2_NUM91_OUT, XNOR_1_2_AND2_NUM91_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM91 (.ZN (XNOR_1_1_AND2_NUM91_OUT), .A1 (N66), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM91 (.ZN (XNOR_1_2_AND2_NUM91_OUT), .A1 (GND), .A2 (N319));
      NOR2_X1 XNOR_1_3_AND2_NUM91 (.ZN (N586), .A1 (XNOR_1_1_AND2_NUM91_OUT), .A2 (XNOR_1_2_AND2_NUM91_OUT));
      wire XNOR_1_1_BUFF1_NUM92_OUT;
      NOR2_X1 XNOR_1_1_BUFF1_NUM92 (.ZN (XNOR_1_1_BUFF1_NUM92_OUT), .A1 (N239), .A2 (GND));
      NOR2_X1 XNOR_1_2_BUFF1_NUM92 (.ZN (N589), .A1 (XNOR_1_1_BUFF1_NUM92_OUT), .A2 (GND));
      wire XNOR_1_1_AND3_NUM93_OUT, XNOR_1_2_AND3_NUM93_OUT, XNOR_1_3_AND3_NUM93_OUT;
      NOR2_X1 XNOR_1_1_AND3_NUM93 (.ZN (XNOR_1_1_AND3_NUM93_OUT), .A1 (N49), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND3_NUM93 (.ZN (XNOR_1_2_AND3_NUM93_OUT), .A1 (GND), .A2 (N253));
      NOR2_X1 XNOR_1_3_AND3_NUM93 (.ZN (XNOR_1_3_AND3_NUM93_OUT), .A1 (XNOR_1_1_AND3_NUM93_OUT), .A2 (XNOR_1_2_AND3_NUM93_OUT));

      wire XNOR_2_1_AND3_NUM93_OUT, XNOR_2_2_AND3_NUM93_OUT;
      NOR2_X1 XNOR_2_1_AND3_NUM93 (.ZN (XNOR_2_1_AND3_NUM93_OUT), .A1 (N319), .A2 (GND));
      NOR2_X1 XNOR_2_2_AND3_NUM93 (.ZN (XNOR_2_2_AND3_NUM93_OUT), .A1 (GND), .A2 (XNOR_1_3_AND3_NUM93_OUT));
      NOR2_X1 XNOR_2_3_AND3_NUM93 (.ZN (N592), .A1 (XNOR_2_1_AND3_NUM93_OUT), .A2 (XNOR_2_2_AND3_NUM93_OUT));
      wire XNOR_1_1_BUFF1_NUM94_OUT;
      NOR2_X1 XNOR_1_1_BUFF1_NUM94 (.ZN (XNOR_1_1_BUFF1_NUM94_OUT), .A1 (N247), .A2 (GND));
      NOR2_X1 XNOR_1_2_BUFF1_NUM94 (.ZN (N595), .A1 (XNOR_1_1_BUFF1_NUM94_OUT), .A2 (GND));
      wire XNOR_1_1_BUFF1_NUM95_OUT;
      NOR2_X1 XNOR_1_1_BUFF1_NUM95 (.ZN (XNOR_1_1_BUFF1_NUM95_OUT), .A1 (N239), .A2 (GND));
      NOR2_X1 XNOR_1_2_BUFF1_NUM95 (.ZN (N598), .A1 (XNOR_1_1_BUFF1_NUM95_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM96_OUT, XNOR_1_2_NAND2_NUM96_OUT, XNOR_1_3_NAND2_NUM96_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM96 (.ZN (XNOR_1_1_NAND2_NUM96_OUT), .A1 (N326), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM96 (.ZN (XNOR_1_2_NAND2_NUM96_OUT), .A1 (GND), .A2 (N277));
      NOR2_X1 XNOR_1_3_NAND2_NUM96 (.ZN (XNOR_1_3_NAND2_NUM96_OUT), .A1 (XNOR_1_1_NAND2_NUM96_OUT), .A2 (XNOR_1_2_NAND2_NUM96_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM96 (.ZN (N601), .A1 (XNOR_1_3_NAND2_NUM96_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM97_OUT, XNOR_1_2_NAND2_NUM97_OUT, XNOR_1_3_NAND2_NUM97_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM97 (.ZN (XNOR_1_1_NAND2_NUM97_OUT), .A1 (N326), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM97 (.ZN (XNOR_1_2_NAND2_NUM97_OUT), .A1 (GND), .A2 (N280));
      NOR2_X1 XNOR_1_3_NAND2_NUM97 (.ZN (XNOR_1_3_NAND2_NUM97_OUT), .A1 (XNOR_1_1_NAND2_NUM97_OUT), .A2 (XNOR_1_2_NAND2_NUM97_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM97 (.ZN (N602), .A1 (XNOR_1_3_NAND2_NUM97_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM98_OUT, XNOR_1_2_NAND2_NUM98_OUT, XNOR_1_3_NAND2_NUM98_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM98 (.ZN (XNOR_1_1_NAND2_NUM98_OUT), .A1 (N260), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM98 (.ZN (XNOR_1_2_NAND2_NUM98_OUT), .A1 (GND), .A2 (N72));
      NOR2_X1 XNOR_1_3_NAND2_NUM98 (.ZN (XNOR_1_3_NAND2_NUM98_OUT), .A1 (XNOR_1_1_NAND2_NUM98_OUT), .A2 (XNOR_1_2_NAND2_NUM98_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM98 (.ZN (N603), .A1 (XNOR_1_3_NAND2_NUM98_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM99_OUT, XNOR_1_2_NAND2_NUM99_OUT, XNOR_1_3_NAND2_NUM99_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM99 (.ZN (XNOR_1_1_NAND2_NUM99_OUT), .A1 (N260), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM99 (.ZN (XNOR_1_2_NAND2_NUM99_OUT), .A1 (GND), .A2 (N300));
      NOR2_X1 XNOR_1_3_NAND2_NUM99 (.ZN (XNOR_1_3_NAND2_NUM99_OUT), .A1 (XNOR_1_1_NAND2_NUM99_OUT), .A2 (XNOR_1_2_NAND2_NUM99_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM99 (.ZN (N608), .A1 (XNOR_1_3_NAND2_NUM99_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM100_OUT, XNOR_1_2_NAND2_NUM100_OUT, XNOR_1_3_NAND2_NUM100_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM100 (.ZN (XNOR_1_1_NAND2_NUM100_OUT), .A1 (N256), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM100 (.ZN (XNOR_1_2_NAND2_NUM100_OUT), .A1 (GND), .A2 (N300));
      NOR2_X1 XNOR_1_3_NAND2_NUM100 (.ZN (XNOR_1_3_NAND2_NUM100_OUT), .A1 (XNOR_1_1_NAND2_NUM100_OUT), .A2 (XNOR_1_2_NAND2_NUM100_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM100 (.ZN (N612), .A1 (XNOR_1_3_NAND2_NUM100_OUT), .A2 (GND));
      wire XNOR_1_1_BUFF1_NUM101_OUT;
      NOR2_X1 XNOR_1_1_BUFF1_NUM101 (.ZN (XNOR_1_1_BUFF1_NUM101_OUT), .A1 (N201), .A2 (GND));
      NOR2_X1 XNOR_1_2_BUFF1_NUM101 (.ZN (N616), .A1 (XNOR_1_1_BUFF1_NUM101_OUT), .A2 (GND));
      wire XNOR_1_1_BUFF1_NUM102_OUT;
      NOR2_X1 XNOR_1_1_BUFF1_NUM102 (.ZN (XNOR_1_1_BUFF1_NUM102_OUT), .A1 (N216), .A2 (GND));
      NOR2_X1 XNOR_1_2_BUFF1_NUM102 (.ZN (N619), .A1 (XNOR_1_1_BUFF1_NUM102_OUT), .A2 (GND));
      wire XNOR_1_1_BUFF1_NUM103_OUT;
      NOR2_X1 XNOR_1_1_BUFF1_NUM103 (.ZN (XNOR_1_1_BUFF1_NUM103_OUT), .A1 (N220), .A2 (GND));
      NOR2_X1 XNOR_1_2_BUFF1_NUM103 (.ZN (N622), .A1 (XNOR_1_1_BUFF1_NUM103_OUT), .A2 (GND));
      wire XNOR_1_1_BUFF1_NUM104_OUT;
      NOR2_X1 XNOR_1_1_BUFF1_NUM104 (.ZN (XNOR_1_1_BUFF1_NUM104_OUT), .A1 (N239), .A2 (GND));
      NOR2_X1 XNOR_1_2_BUFF1_NUM104 (.ZN (N625), .A1 (XNOR_1_1_BUFF1_NUM104_OUT), .A2 (GND));
      wire XNOR_1_1_BUFF1_NUM105_OUT;
      NOR2_X1 XNOR_1_1_BUFF1_NUM105 (.ZN (XNOR_1_1_BUFF1_NUM105_OUT), .A1 (N190), .A2 (GND));
      NOR2_X1 XNOR_1_2_BUFF1_NUM105 (.ZN (N628), .A1 (XNOR_1_1_BUFF1_NUM105_OUT), .A2 (GND));
      wire XNOR_1_1_BUFF1_NUM106_OUT;
      NOR2_X1 XNOR_1_1_BUFF1_NUM106 (.ZN (XNOR_1_1_BUFF1_NUM106_OUT), .A1 (N190), .A2 (GND));
      NOR2_X1 XNOR_1_2_BUFF1_NUM106 (.ZN (N631), .A1 (XNOR_1_1_BUFF1_NUM106_OUT), .A2 (GND));
      wire XNOR_1_1_BUFF1_NUM107_OUT;
      NOR2_X1 XNOR_1_1_BUFF1_NUM107 (.ZN (XNOR_1_1_BUFF1_NUM107_OUT), .A1 (N194), .A2 (GND));
      NOR2_X1 XNOR_1_2_BUFF1_NUM107 (.ZN (N634), .A1 (XNOR_1_1_BUFF1_NUM107_OUT), .A2 (GND));
      wire XNOR_1_1_BUFF1_NUM108_OUT;
      NOR2_X1 XNOR_1_1_BUFF1_NUM108 (.ZN (XNOR_1_1_BUFF1_NUM108_OUT), .A1 (N229), .A2 (GND));
      NOR2_X1 XNOR_1_2_BUFF1_NUM108 (.ZN (N637), .A1 (XNOR_1_1_BUFF1_NUM108_OUT), .A2 (GND));
      wire XNOR_1_1_BUFF1_NUM109_OUT;
      NOR2_X1 XNOR_1_1_BUFF1_NUM109 (.ZN (XNOR_1_1_BUFF1_NUM109_OUT), .A1 (N197), .A2 (GND));
      NOR2_X1 XNOR_1_2_BUFF1_NUM109 (.ZN (N640), .A1 (XNOR_1_1_BUFF1_NUM109_OUT), .A2 (GND));
      wire XNOR_1_1_AND3_NUM110_OUT, XNOR_1_2_AND3_NUM110_OUT, XNOR_1_3_AND3_NUM110_OUT;
      NOR2_X1 XNOR_1_1_AND3_NUM110 (.ZN (XNOR_1_1_AND3_NUM110_OUT), .A1 (N56), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND3_NUM110 (.ZN (XNOR_1_2_AND3_NUM110_OUT), .A1 (GND), .A2 (N257));
      NOR2_X1 XNOR_1_3_AND3_NUM110 (.ZN (XNOR_1_3_AND3_NUM110_OUT), .A1 (XNOR_1_1_AND3_NUM110_OUT), .A2 (XNOR_1_2_AND3_NUM110_OUT));

      wire XNOR_2_1_AND3_NUM110_OUT, XNOR_2_2_AND3_NUM110_OUT;
      NOR2_X1 XNOR_2_1_AND3_NUM110 (.ZN (XNOR_2_1_AND3_NUM110_OUT), .A1 (N319), .A2 (GND));
      NOR2_X1 XNOR_2_2_AND3_NUM110 (.ZN (XNOR_2_2_AND3_NUM110_OUT), .A1 (GND), .A2 (XNOR_1_3_AND3_NUM110_OUT));
      NOR2_X1 XNOR_2_3_AND3_NUM110 (.ZN (N643), .A1 (XNOR_2_1_AND3_NUM110_OUT), .A2 (XNOR_2_2_AND3_NUM110_OUT));
      wire XNOR_1_1_BUFF1_NUM111_OUT;
      NOR2_X1 XNOR_1_1_BUFF1_NUM111 (.ZN (XNOR_1_1_BUFF1_NUM111_OUT), .A1 (N232), .A2 (GND));
      NOR2_X1 XNOR_1_2_BUFF1_NUM111 (.ZN (N646), .A1 (XNOR_1_1_BUFF1_NUM111_OUT), .A2 (GND));
      wire XNOR_1_1_BUFF1_NUM112_OUT;
      NOR2_X1 XNOR_1_1_BUFF1_NUM112 (.ZN (XNOR_1_1_BUFF1_NUM112_OUT), .A1 (N201), .A2 (GND));
      NOR2_X1 XNOR_1_2_BUFF1_NUM112 (.ZN (N649), .A1 (XNOR_1_1_BUFF1_NUM112_OUT), .A2 (GND));
      wire XNOR_1_1_BUFF1_NUM113_OUT;
      NOR2_X1 XNOR_1_1_BUFF1_NUM113 (.ZN (XNOR_1_1_BUFF1_NUM113_OUT), .A1 (N235), .A2 (GND));
      NOR2_X1 XNOR_1_2_BUFF1_NUM113 (.ZN (N652), .A1 (XNOR_1_1_BUFF1_NUM113_OUT), .A2 (GND));
      wire XNOR_1_1_AND3_NUM114_OUT, XNOR_1_2_AND3_NUM114_OUT, XNOR_1_3_AND3_NUM114_OUT;
      NOR2_X1 XNOR_1_1_AND3_NUM114 (.ZN (XNOR_1_1_AND3_NUM114_OUT), .A1 (N60), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND3_NUM114 (.ZN (XNOR_1_2_AND3_NUM114_OUT), .A1 (GND), .A2 (N257));
      NOR2_X1 XNOR_1_3_AND3_NUM114 (.ZN (XNOR_1_3_AND3_NUM114_OUT), .A1 (XNOR_1_1_AND3_NUM114_OUT), .A2 (XNOR_1_2_AND3_NUM114_OUT));

      wire XNOR_2_1_AND3_NUM114_OUT, XNOR_2_2_AND3_NUM114_OUT;
      NOR2_X1 XNOR_2_1_AND3_NUM114 (.ZN (XNOR_2_1_AND3_NUM114_OUT), .A1 (N319), .A2 (GND));
      NOR2_X1 XNOR_2_2_AND3_NUM114 (.ZN (XNOR_2_2_AND3_NUM114_OUT), .A1 (GND), .A2 (XNOR_1_3_AND3_NUM114_OUT));
      NOR2_X1 XNOR_2_3_AND3_NUM114 (.ZN (N655), .A1 (XNOR_2_1_AND3_NUM114_OUT), .A2 (XNOR_2_2_AND3_NUM114_OUT));
      wire XNOR_1_1_BUFF1_NUM115_OUT;
      NOR2_X1 XNOR_1_1_BUFF1_NUM115 (.ZN (XNOR_1_1_BUFF1_NUM115_OUT), .A1 (N263), .A2 (GND));
      NOR2_X1 XNOR_1_2_BUFF1_NUM115 (.ZN (N658), .A1 (XNOR_1_1_BUFF1_NUM115_OUT), .A2 (GND));
      wire XNOR_1_1_BUFF1_NUM116_OUT;
      NOR2_X1 XNOR_1_1_BUFF1_NUM116 (.ZN (XNOR_1_1_BUFF1_NUM116_OUT), .A1 (N263), .A2 (GND));
      NOR2_X1 XNOR_1_2_BUFF1_NUM116 (.ZN (N661), .A1 (XNOR_1_1_BUFF1_NUM116_OUT), .A2 (GND));
      wire XNOR_1_1_BUFF1_NUM117_OUT;
      NOR2_X1 XNOR_1_1_BUFF1_NUM117 (.ZN (XNOR_1_1_BUFF1_NUM117_OUT), .A1 (N266), .A2 (GND));
      NOR2_X1 XNOR_1_2_BUFF1_NUM117 (.ZN (N664), .A1 (XNOR_1_1_BUFF1_NUM117_OUT), .A2 (GND));
      wire XNOR_1_1_BUFF1_NUM118_OUT;
      NOR2_X1 XNOR_1_1_BUFF1_NUM118 (.ZN (XNOR_1_1_BUFF1_NUM118_OUT), .A1 (N266), .A2 (GND));
      NOR2_X1 XNOR_1_2_BUFF1_NUM118 (.ZN (N667), .A1 (XNOR_1_1_BUFF1_NUM118_OUT), .A2 (GND));
      wire XNOR_1_1_BUFF1_NUM119_OUT;
      NOR2_X1 XNOR_1_1_BUFF1_NUM119 (.ZN (XNOR_1_1_BUFF1_NUM119_OUT), .A1 (N269), .A2 (GND));
      NOR2_X1 XNOR_1_2_BUFF1_NUM119 (.ZN (N670), .A1 (XNOR_1_1_BUFF1_NUM119_OUT), .A2 (GND));
      wire XNOR_1_1_BUFF1_NUM120_OUT;
      NOR2_X1 XNOR_1_1_BUFF1_NUM120 (.ZN (XNOR_1_1_BUFF1_NUM120_OUT), .A1 (N269), .A2 (GND));
      NOR2_X1 XNOR_1_2_BUFF1_NUM120 (.ZN (N673), .A1 (XNOR_1_1_BUFF1_NUM120_OUT), .A2 (GND));
      wire XNOR_1_1_BUFF1_NUM121_OUT;
      NOR2_X1 XNOR_1_1_BUFF1_NUM121 (.ZN (XNOR_1_1_BUFF1_NUM121_OUT), .A1 (N272), .A2 (GND));
      NOR2_X1 XNOR_1_2_BUFF1_NUM121 (.ZN (N676), .A1 (XNOR_1_1_BUFF1_NUM121_OUT), .A2 (GND));
      wire XNOR_1_1_BUFF1_NUM122_OUT;
      NOR2_X1 XNOR_1_1_BUFF1_NUM122 (.ZN (XNOR_1_1_BUFF1_NUM122_OUT), .A1 (N272), .A2 (GND));
      NOR2_X1 XNOR_1_2_BUFF1_NUM122 (.ZN (N679), .A1 (XNOR_1_1_BUFF1_NUM122_OUT), .A2 (GND));
      wire XNOR_1_1_AND2_NUM123_OUT, XNOR_1_2_AND2_NUM123_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM123 (.ZN (XNOR_1_1_AND2_NUM123_OUT), .A1 (N251), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM123 (.ZN (XNOR_1_2_AND2_NUM123_OUT), .A1 (GND), .A2 (N316));
      NOR2_X1 XNOR_1_3_AND2_NUM123 (.ZN (N682), .A1 (XNOR_1_1_AND2_NUM123_OUT), .A2 (XNOR_1_2_AND2_NUM123_OUT));
      wire XNOR_1_1_AND2_NUM124_OUT, XNOR_1_2_AND2_NUM124_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM124 (.ZN (XNOR_1_1_AND2_NUM124_OUT), .A1 (N252), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM124 (.ZN (XNOR_1_2_AND2_NUM124_OUT), .A1 (GND), .A2 (N316));
      NOR2_X1 XNOR_1_3_AND2_NUM124 (.ZN (N685), .A1 (XNOR_1_1_AND2_NUM124_OUT), .A2 (XNOR_1_2_AND2_NUM124_OUT));
      wire XNOR_1_1_BUFF1_NUM125_OUT;
      NOR2_X1 XNOR_1_1_BUFF1_NUM125 (.ZN (XNOR_1_1_BUFF1_NUM125_OUT), .A1 (N197), .A2 (GND));
      NOR2_X1 XNOR_1_2_BUFF1_NUM125 (.ZN (N688), .A1 (XNOR_1_1_BUFF1_NUM125_OUT), .A2 (GND));
      wire XNOR_1_1_BUFF1_NUM126_OUT;
      NOR2_X1 XNOR_1_1_BUFF1_NUM126 (.ZN (XNOR_1_1_BUFF1_NUM126_OUT), .A1 (N197), .A2 (GND));
      NOR2_X1 XNOR_1_2_BUFF1_NUM126 (.ZN (N691), .A1 (XNOR_1_1_BUFF1_NUM126_OUT), .A2 (GND));
      wire XNOR_1_1_BUFF1_NUM127_OUT;
      NOR2_X1 XNOR_1_1_BUFF1_NUM127 (.ZN (XNOR_1_1_BUFF1_NUM127_OUT), .A1 (N212), .A2 (GND));
      NOR2_X1 XNOR_1_2_BUFF1_NUM127 (.ZN (N694), .A1 (XNOR_1_1_BUFF1_NUM127_OUT), .A2 (GND));
      wire XNOR_1_1_BUFF1_NUM128_OUT;
      NOR2_X1 XNOR_1_1_BUFF1_NUM128 (.ZN (XNOR_1_1_BUFF1_NUM128_OUT), .A1 (N212), .A2 (GND));
      NOR2_X1 XNOR_1_2_BUFF1_NUM128 (.ZN (N697), .A1 (XNOR_1_1_BUFF1_NUM128_OUT), .A2 (GND));
      wire XNOR_1_1_BUFF1_NUM129_OUT;
      NOR2_X1 XNOR_1_1_BUFF1_NUM129 (.ZN (XNOR_1_1_BUFF1_NUM129_OUT), .A1 (N247), .A2 (GND));
      NOR2_X1 XNOR_1_2_BUFF1_NUM129 (.ZN (N700), .A1 (XNOR_1_1_BUFF1_NUM129_OUT), .A2 (GND));
      wire XNOR_1_1_BUFF1_NUM130_OUT;
      NOR2_X1 XNOR_1_1_BUFF1_NUM130 (.ZN (XNOR_1_1_BUFF1_NUM130_OUT), .A1 (N247), .A2 (GND));
      NOR2_X1 XNOR_1_2_BUFF1_NUM130 (.ZN (N703), .A1 (XNOR_1_1_BUFF1_NUM130_OUT), .A2 (GND));
      wire XNOR_1_1_BUFF1_NUM131_OUT;
      NOR2_X1 XNOR_1_1_BUFF1_NUM131 (.ZN (XNOR_1_1_BUFF1_NUM131_OUT), .A1 (N235), .A2 (GND));
      NOR2_X1 XNOR_1_2_BUFF1_NUM131 (.ZN (N706), .A1 (XNOR_1_1_BUFF1_NUM131_OUT), .A2 (GND));
      wire XNOR_1_1_BUFF1_NUM132_OUT;
      NOR2_X1 XNOR_1_1_BUFF1_NUM132 (.ZN (XNOR_1_1_BUFF1_NUM132_OUT), .A1 (N235), .A2 (GND));
      NOR2_X1 XNOR_1_2_BUFF1_NUM132 (.ZN (N709), .A1 (XNOR_1_1_BUFF1_NUM132_OUT), .A2 (GND));
      wire XNOR_1_1_BUFF1_NUM133_OUT;
      NOR2_X1 XNOR_1_1_BUFF1_NUM133 (.ZN (XNOR_1_1_BUFF1_NUM133_OUT), .A1 (N201), .A2 (GND));
      NOR2_X1 XNOR_1_2_BUFF1_NUM133 (.ZN (N712), .A1 (XNOR_1_1_BUFF1_NUM133_OUT), .A2 (GND));
      wire XNOR_1_1_BUFF1_NUM134_OUT;
      NOR2_X1 XNOR_1_1_BUFF1_NUM134 (.ZN (XNOR_1_1_BUFF1_NUM134_OUT), .A1 (N201), .A2 (GND));
      NOR2_X1 XNOR_1_2_BUFF1_NUM134 (.ZN (N715), .A1 (XNOR_1_1_BUFF1_NUM134_OUT), .A2 (GND));
      wire XNOR_1_1_BUFF1_NUM135_OUT;
      NOR2_X1 XNOR_1_1_BUFF1_NUM135 (.ZN (XNOR_1_1_BUFF1_NUM135_OUT), .A1 (N206), .A2 (GND));
      NOR2_X1 XNOR_1_2_BUFF1_NUM135 (.ZN (N718), .A1 (XNOR_1_1_BUFF1_NUM135_OUT), .A2 (GND));
      wire XNOR_1_1_BUFF1_NUM136_OUT;
      NOR2_X1 XNOR_1_1_BUFF1_NUM136 (.ZN (XNOR_1_1_BUFF1_NUM136_OUT), .A1 (N216), .A2 (GND));
      NOR2_X1 XNOR_1_2_BUFF1_NUM136 (.ZN (N721), .A1 (XNOR_1_1_BUFF1_NUM136_OUT), .A2 (GND));
      wire XNOR_1_1_AND3_NUM137_OUT, XNOR_1_2_AND3_NUM137_OUT, XNOR_1_3_AND3_NUM137_OUT;
      NOR2_X1 XNOR_1_1_AND3_NUM137 (.ZN (XNOR_1_1_AND3_NUM137_OUT), .A1 (N53), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND3_NUM137 (.ZN (XNOR_1_2_AND3_NUM137_OUT), .A1 (GND), .A2 (N253));
      NOR2_X1 XNOR_1_3_AND3_NUM137 (.ZN (XNOR_1_3_AND3_NUM137_OUT), .A1 (XNOR_1_1_AND3_NUM137_OUT), .A2 (XNOR_1_2_AND3_NUM137_OUT));

      wire XNOR_2_1_AND3_NUM137_OUT, XNOR_2_2_AND3_NUM137_OUT;
      NOR2_X1 XNOR_2_1_AND3_NUM137 (.ZN (XNOR_2_1_AND3_NUM137_OUT), .A1 (N319), .A2 (GND));
      NOR2_X1 XNOR_2_2_AND3_NUM137 (.ZN (XNOR_2_2_AND3_NUM137_OUT), .A1 (GND), .A2 (XNOR_1_3_AND3_NUM137_OUT));
      NOR2_X1 XNOR_2_3_AND3_NUM137 (.ZN (N724), .A1 (XNOR_2_1_AND3_NUM137_OUT), .A2 (XNOR_2_2_AND3_NUM137_OUT));
      wire XNOR_1_1_BUFF1_NUM138_OUT;
      NOR2_X1 XNOR_1_1_BUFF1_NUM138 (.ZN (XNOR_1_1_BUFF1_NUM138_OUT), .A1 (N243), .A2 (GND));
      NOR2_X1 XNOR_1_2_BUFF1_NUM138 (.ZN (N727), .A1 (XNOR_1_1_BUFF1_NUM138_OUT), .A2 (GND));
      wire XNOR_1_1_BUFF1_NUM139_OUT;
      NOR2_X1 XNOR_1_1_BUFF1_NUM139 (.ZN (XNOR_1_1_BUFF1_NUM139_OUT), .A1 (N220), .A2 (GND));
      NOR2_X1 XNOR_1_2_BUFF1_NUM139 (.ZN (N730), .A1 (XNOR_1_1_BUFF1_NUM139_OUT), .A2 (GND));
      wire XNOR_1_1_BUFF1_NUM140_OUT;
      NOR2_X1 XNOR_1_1_BUFF1_NUM140 (.ZN (XNOR_1_1_BUFF1_NUM140_OUT), .A1 (N220), .A2 (GND));
      NOR2_X1 XNOR_1_2_BUFF1_NUM140 (.ZN (N733), .A1 (XNOR_1_1_BUFF1_NUM140_OUT), .A2 (GND));
      wire XNOR_1_1_BUFF1_NUM141_OUT;
      NOR2_X1 XNOR_1_1_BUFF1_NUM141 (.ZN (XNOR_1_1_BUFF1_NUM141_OUT), .A1 (N209), .A2 (GND));
      NOR2_X1 XNOR_1_2_BUFF1_NUM141 (.ZN (N736), .A1 (XNOR_1_1_BUFF1_NUM141_OUT), .A2 (GND));
      wire XNOR_1_1_BUFF1_NUM142_OUT;
      NOR2_X1 XNOR_1_1_BUFF1_NUM142 (.ZN (XNOR_1_1_BUFF1_NUM142_OUT), .A1 (N216), .A2 (GND));
      NOR2_X1 XNOR_1_2_BUFF1_NUM142 (.ZN (N739), .A1 (XNOR_1_1_BUFF1_NUM142_OUT), .A2 (GND));
      wire XNOR_1_1_BUFF1_NUM143_OUT;
      NOR2_X1 XNOR_1_1_BUFF1_NUM143 (.ZN (XNOR_1_1_BUFF1_NUM143_OUT), .A1 (N225), .A2 (GND));
      NOR2_X1 XNOR_1_2_BUFF1_NUM143 (.ZN (N742), .A1 (XNOR_1_1_BUFF1_NUM143_OUT), .A2 (GND));
      wire XNOR_1_1_BUFF1_NUM144_OUT;
      NOR2_X1 XNOR_1_1_BUFF1_NUM144 (.ZN (XNOR_1_1_BUFF1_NUM144_OUT), .A1 (N243), .A2 (GND));
      NOR2_X1 XNOR_1_2_BUFF1_NUM144 (.ZN (N745), .A1 (XNOR_1_1_BUFF1_NUM144_OUT), .A2 (GND));
      wire XNOR_1_1_BUFF1_NUM145_OUT;
      NOR2_X1 XNOR_1_1_BUFF1_NUM145 (.ZN (XNOR_1_1_BUFF1_NUM145_OUT), .A1 (N212), .A2 (GND));
      NOR2_X1 XNOR_1_2_BUFF1_NUM145 (.ZN (N748), .A1 (XNOR_1_1_BUFF1_NUM145_OUT), .A2 (GND));
      wire XNOR_1_1_BUFF1_NUM146_OUT;
      NOR2_X1 XNOR_1_1_BUFF1_NUM146 (.ZN (XNOR_1_1_BUFF1_NUM146_OUT), .A1 (N225), .A2 (GND));
      NOR2_X1 XNOR_1_2_BUFF1_NUM146 (.ZN (N751), .A1 (XNOR_1_1_BUFF1_NUM146_OUT), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM147 (.ZN (N886), .A1 (N682), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM148 (.ZN (N887), .A1 (N685), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM149 (.ZN (N888), .A1 (N616), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM150 (.ZN (N889), .A1 (N619), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM151 (.ZN (N890), .A1 (N622), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM152 (.ZN (N891), .A1 (N625), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM153 (.ZN (N892), .A1 (N631), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM154 (.ZN (N893), .A1 (N643), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM155 (.ZN (N894), .A1 (N649), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM156 (.ZN (N895), .A1 (N652), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM157 (.ZN (N896), .A1 (N655), .A2 (GND));
      wire XNOR_1_1_AND2_NUM158_OUT, XNOR_1_2_AND2_NUM158_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM158 (.ZN (XNOR_1_1_AND2_NUM158_OUT), .A1 (N49), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM158 (.ZN (XNOR_1_2_AND2_NUM158_OUT), .A1 (GND), .A2 (N612));
      NOR2_X1 XNOR_1_3_AND2_NUM158 (.ZN (N897), .A1 (XNOR_1_1_AND2_NUM158_OUT), .A2 (XNOR_1_2_AND2_NUM158_OUT));
      wire XNOR_1_1_AND2_NUM159_OUT, XNOR_1_2_AND2_NUM159_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM159 (.ZN (XNOR_1_1_AND2_NUM159_OUT), .A1 (N56), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM159 (.ZN (XNOR_1_2_AND2_NUM159_OUT), .A1 (GND), .A2 (N608));
      NOR2_X1 XNOR_1_3_AND2_NUM159 (.ZN (N898), .A1 (XNOR_1_1_AND2_NUM159_OUT), .A2 (XNOR_1_2_AND2_NUM159_OUT));
      wire XNOR_1_1_NAND2_NUM160_OUT, XNOR_1_2_NAND2_NUM160_OUT, XNOR_1_3_NAND2_NUM160_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM160 (.ZN (XNOR_1_1_NAND2_NUM160_OUT), .A1 (N53), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM160 (.ZN (XNOR_1_2_NAND2_NUM160_OUT), .A1 (GND), .A2 (N612));
      NOR2_X1 XNOR_1_3_NAND2_NUM160 (.ZN (XNOR_1_3_NAND2_NUM160_OUT), .A1 (XNOR_1_1_NAND2_NUM160_OUT), .A2 (XNOR_1_2_NAND2_NUM160_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM160 (.ZN (N899), .A1 (XNOR_1_3_NAND2_NUM160_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM161_OUT, XNOR_1_2_NAND2_NUM161_OUT, XNOR_1_3_NAND2_NUM161_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM161 (.ZN (XNOR_1_1_NAND2_NUM161_OUT), .A1 (N60), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM161 (.ZN (XNOR_1_2_NAND2_NUM161_OUT), .A1 (GND), .A2 (N608));
      NOR2_X1 XNOR_1_3_NAND2_NUM161 (.ZN (XNOR_1_3_NAND2_NUM161_OUT), .A1 (XNOR_1_1_NAND2_NUM161_OUT), .A2 (XNOR_1_2_NAND2_NUM161_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM161 (.ZN (N903), .A1 (XNOR_1_3_NAND2_NUM161_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM162_OUT, XNOR_1_2_NAND2_NUM162_OUT, XNOR_1_3_NAND2_NUM162_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM162 (.ZN (XNOR_1_1_NAND2_NUM162_OUT), .A1 (N49), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM162 (.ZN (XNOR_1_2_NAND2_NUM162_OUT), .A1 (GND), .A2 (N612));
      NOR2_X1 XNOR_1_3_NAND2_NUM162 (.ZN (XNOR_1_3_NAND2_NUM162_OUT), .A1 (XNOR_1_1_NAND2_NUM162_OUT), .A2 (XNOR_1_2_NAND2_NUM162_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM162 (.ZN (N907), .A1 (XNOR_1_3_NAND2_NUM162_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM163_OUT, XNOR_1_2_NAND2_NUM163_OUT, XNOR_1_3_NAND2_NUM163_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM163 (.ZN (XNOR_1_1_NAND2_NUM163_OUT), .A1 (N56), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM163 (.ZN (XNOR_1_2_NAND2_NUM163_OUT), .A1 (GND), .A2 (N608));
      NOR2_X1 XNOR_1_3_NAND2_NUM163 (.ZN (XNOR_1_3_NAND2_NUM163_OUT), .A1 (XNOR_1_1_NAND2_NUM163_OUT), .A2 (XNOR_1_2_NAND2_NUM163_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM163 (.ZN (N910), .A1 (XNOR_1_3_NAND2_NUM163_OUT), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM164 (.ZN (N913), .A1 (N661), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM165 (.ZN (N914), .A1 (N658), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM166 (.ZN (N915), .A1 (N667), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM167 (.ZN (N916), .A1 (N664), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM168 (.ZN (N917), .A1 (N673), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM169 (.ZN (N918), .A1 (N670), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM170 (.ZN (N919), .A1 (N679), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM171 (.ZN (N920), .A1 (N676), .A2 (GND));
      wire XNOR_1_1_NAND4_NUM172_OUT, XNOR_1_2_NAND4_NUM172_OUT, XNOR_1_3_NAND4_NUM172_OUT;
      NOR2_X1 XNOR_1_1_NAND4_NUM172 (.ZN (XNOR_1_1_NAND4_NUM172_OUT), .A1 (N277), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND4_NUM172 (.ZN (XNOR_1_2_NAND4_NUM172_OUT), .A1 (GND), .A2 (N297));
      NOR2_X1 XNOR_1_3_NAND4_NUM172 (.ZN (XNOR_1_3_NAND4_NUM172_OUT), .A1 (XNOR_1_1_NAND4_NUM172_OUT), .A2 (XNOR_1_2_NAND4_NUM172_OUT));

      wire XNOR_2_1_NAND4_NUM172_OUT, XNOR_2_2_NAND4_NUM172_OUT, XNOR_2_3_NAND4_NUM172_OUT;
      NOR2_X1 XNOR_2_1_NAND4_NUM172 (.ZN (XNOR_2_1_NAND4_NUM172_OUT), .A1 (N326), .A2 (GND));
      NOR2_X1 XNOR_2_2_NAND4_NUM172 (.ZN (XNOR_2_2_NAND4_NUM172_OUT), .A1 (GND), .A2 (N603));
      NOR2_X1 XNOR_2_3_NAND4_NUM172 (.ZN (XNOR_2_3_NAND4_NUM172_OUT), .A1 (XNOR_2_1_NAND4_NUM172_OUT), .A2 (XNOR_2_2_NAND4_NUM172_OUT));

      wire XNOR_3_1_NAND4_NUM172_OUT, XNOR_3_2_NAND4_NUM172_OUT, XNOR_3_3_NAND4_NUM172_OUT;
      NOR2_X1 XNOR_3_1_NAND4_NUM172 (.ZN (XNOR_3_1_NAND4_NUM172_OUT), .A1 (XNOR_1_3_NAND4_NUM172_OUT), .A2 (GND));
      NOR2_X1 XNOR_3_2_NAND4_NUM172 (.ZN (XNOR_3_2_NAND4_NUM172_OUT), .A1 (GND), .A2 (XNOR_2_3_NAND4_NUM172_OUT));
      NOR2_X1 XNOR_3_3_NAND4_NUM172 (.ZN (XNOR_3_3_NAND4_NUM172_OUT), .A1 (XNOR_3_1_NAND4_NUM172_OUT), .A2 (XNOR_3_2_NAND4_NUM172_OUT));

      NOR2_X1 XNOR_4_1_NAND4_NUM172 (.ZN (N921), .A1 (XNOR_3_3_NAND4_NUM172_OUT), .A2 (GND));
      wire XNOR_1_1_NAND4_NUM173_OUT, XNOR_1_2_NAND4_NUM173_OUT, XNOR_1_3_NAND4_NUM173_OUT;
      NOR2_X1 XNOR_1_1_NAND4_NUM173 (.ZN (XNOR_1_1_NAND4_NUM173_OUT), .A1 (N280), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND4_NUM173 (.ZN (XNOR_1_2_NAND4_NUM173_OUT), .A1 (GND), .A2 (N297));
      NOR2_X1 XNOR_1_3_NAND4_NUM173 (.ZN (XNOR_1_3_NAND4_NUM173_OUT), .A1 (XNOR_1_1_NAND4_NUM173_OUT), .A2 (XNOR_1_2_NAND4_NUM173_OUT));

      wire XNOR_2_1_NAND4_NUM173_OUT, XNOR_2_2_NAND4_NUM173_OUT, XNOR_2_3_NAND4_NUM173_OUT;
      NOR2_X1 XNOR_2_1_NAND4_NUM173 (.ZN (XNOR_2_1_NAND4_NUM173_OUT), .A1 (N326), .A2 (GND));
      NOR2_X1 XNOR_2_2_NAND4_NUM173 (.ZN (XNOR_2_2_NAND4_NUM173_OUT), .A1 (GND), .A2 (N603));
      NOR2_X1 XNOR_2_3_NAND4_NUM173 (.ZN (XNOR_2_3_NAND4_NUM173_OUT), .A1 (XNOR_2_1_NAND4_NUM173_OUT), .A2 (XNOR_2_2_NAND4_NUM173_OUT));

      wire XNOR_3_1_NAND4_NUM173_OUT, XNOR_3_2_NAND4_NUM173_OUT, XNOR_3_3_NAND4_NUM173_OUT;
      NOR2_X1 XNOR_3_1_NAND4_NUM173 (.ZN (XNOR_3_1_NAND4_NUM173_OUT), .A1 (XNOR_1_3_NAND4_NUM173_OUT), .A2 (GND));
      NOR2_X1 XNOR_3_2_NAND4_NUM173 (.ZN (XNOR_3_2_NAND4_NUM173_OUT), .A1 (GND), .A2 (XNOR_2_3_NAND4_NUM173_OUT));
      NOR2_X1 XNOR_3_3_NAND4_NUM173 (.ZN (XNOR_3_3_NAND4_NUM173_OUT), .A1 (XNOR_3_1_NAND4_NUM173_OUT), .A2 (XNOR_3_2_NAND4_NUM173_OUT));

      NOR2_X1 XNOR_4_1_NAND4_NUM173 (.ZN (N922), .A1 (XNOR_3_3_NAND4_NUM173_OUT), .A2 (GND));
      wire XNOR_1_1_NAND3_NUM174_OUT, XNOR_1_2_NAND3_NUM174_OUT, XNOR_1_3_NAND3_NUM174_OUT;
      NOR2_X1 XNOR_1_1_NAND3_NUM174 (.ZN (XNOR_1_1_NAND3_NUM174_OUT), .A1 (N303), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND3_NUM174 (.ZN (XNOR_1_2_NAND3_NUM174_OUT), .A1 (GND), .A2 (N338));
      NOR2_X1 XNOR_1_3_NAND3_NUM174 (.ZN (XNOR_1_3_NAND3_NUM174_OUT), .A1 (XNOR_1_1_NAND3_NUM174_OUT), .A2 (XNOR_1_2_NAND3_NUM174_OUT));

      wire XNOR_2_1_NAND3_NUM174_OUT, XNOR_2_2_NAND3_NUM174_OUT, XNOR_2_3_NAND3_NUM174_OUT;
      NOR2_X1 XNOR_2_1_NAND3_NUM174 (.ZN (XNOR_2_1_NAND3_NUM174_OUT), .A1 (N603), .A2 (GND));
      NOR2_X1 XNOR_2_2_NAND3_NUM174 (.ZN (XNOR_2_2_NAND3_NUM174_OUT), .A1 (GND), .A2 (XNOR_1_3_NAND3_NUM174_OUT));
      NOR2_X1 XNOR_2_3_NAND3_NUM174 (.ZN (XNOR_2_3_NAND3_NUM174_OUT), .A1 (XNOR_2_1_NAND3_NUM174_OUT), .A2 (XNOR_2_2_NAND3_NUM174_OUT));

      NOR2_X1 XNOR_3_1_NAND3_NUM174 (.ZN (N923), .A1 (XNOR_2_3_NAND3_NUM174_OUT), .A2 (GND));
      wire XNOR_1_1_AND3_NUM175_OUT, XNOR_1_2_AND3_NUM175_OUT, XNOR_1_3_AND3_NUM175_OUT;
      NOR2_X1 XNOR_1_1_AND3_NUM175 (.ZN (XNOR_1_1_AND3_NUM175_OUT), .A1 (N303), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND3_NUM175 (.ZN (XNOR_1_2_AND3_NUM175_OUT), .A1 (GND), .A2 (N338));
      NOR2_X1 XNOR_1_3_AND3_NUM175 (.ZN (XNOR_1_3_AND3_NUM175_OUT), .A1 (XNOR_1_1_AND3_NUM175_OUT), .A2 (XNOR_1_2_AND3_NUM175_OUT));

      wire XNOR_2_1_AND3_NUM175_OUT, XNOR_2_2_AND3_NUM175_OUT;
      NOR2_X1 XNOR_2_1_AND3_NUM175 (.ZN (XNOR_2_1_AND3_NUM175_OUT), .A1 (N603), .A2 (GND));
      NOR2_X1 XNOR_2_2_AND3_NUM175 (.ZN (XNOR_2_2_AND3_NUM175_OUT), .A1 (GND), .A2 (XNOR_1_3_AND3_NUM175_OUT));
      NOR2_X1 XNOR_2_3_AND3_NUM175 (.ZN (N926), .A1 (XNOR_2_1_AND3_NUM175_OUT), .A2 (XNOR_2_2_AND3_NUM175_OUT));
      wire XNOR_1_1_BUFF1_NUM176_OUT;
      NOR2_X1 XNOR_1_1_BUFF1_NUM176 (.ZN (XNOR_1_1_BUFF1_NUM176_OUT), .A1 (N556), .A2 (GND));
      NOR2_X1 XNOR_1_2_BUFF1_NUM176 (.ZN (N935), .A1 (XNOR_1_1_BUFF1_NUM176_OUT), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM177 (.ZN (N938), .A1 (N688), .A2 (GND));
      wire XNOR_1_1_BUFF1_NUM178_OUT;
      NOR2_X1 XNOR_1_1_BUFF1_NUM178 (.ZN (XNOR_1_1_BUFF1_NUM178_OUT), .A1 (N556), .A2 (GND));
      NOR2_X1 XNOR_1_2_BUFF1_NUM178 (.ZN (N939), .A1 (XNOR_1_1_BUFF1_NUM178_OUT), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM179 (.ZN (N942), .A1 (N691), .A2 (GND));
      wire XNOR_1_1_BUFF1_NUM180_OUT;
      NOR2_X1 XNOR_1_1_BUFF1_NUM180 (.ZN (XNOR_1_1_BUFF1_NUM180_OUT), .A1 (N562), .A2 (GND));
      NOR2_X1 XNOR_1_2_BUFF1_NUM180 (.ZN (N943), .A1 (XNOR_1_1_BUFF1_NUM180_OUT), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM181 (.ZN (N946), .A1 (N694), .A2 (GND));
      wire XNOR_1_1_BUFF1_NUM182_OUT;
      NOR2_X1 XNOR_1_1_BUFF1_NUM182 (.ZN (XNOR_1_1_BUFF1_NUM182_OUT), .A1 (N562), .A2 (GND));
      NOR2_X1 XNOR_1_2_BUFF1_NUM182 (.ZN (N947), .A1 (XNOR_1_1_BUFF1_NUM182_OUT), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM183 (.ZN (N950), .A1 (N697), .A2 (GND));
      wire XNOR_1_1_BUFF1_NUM184_OUT;
      NOR2_X1 XNOR_1_1_BUFF1_NUM184 (.ZN (XNOR_1_1_BUFF1_NUM184_OUT), .A1 (N568), .A2 (GND));
      NOR2_X1 XNOR_1_2_BUFF1_NUM184 (.ZN (N951), .A1 (XNOR_1_1_BUFF1_NUM184_OUT), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM185 (.ZN (N954), .A1 (N700), .A2 (GND));
      wire XNOR_1_1_BUFF1_NUM186_OUT;
      NOR2_X1 XNOR_1_1_BUFF1_NUM186 (.ZN (XNOR_1_1_BUFF1_NUM186_OUT), .A1 (N568), .A2 (GND));
      NOR2_X1 XNOR_1_2_BUFF1_NUM186 (.ZN (N955), .A1 (XNOR_1_1_BUFF1_NUM186_OUT), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM187 (.ZN (N958), .A1 (N703), .A2 (GND));
      wire XNOR_1_1_BUFF1_NUM188_OUT;
      NOR2_X1 XNOR_1_1_BUFF1_NUM188 (.ZN (XNOR_1_1_BUFF1_NUM188_OUT), .A1 (N574), .A2 (GND));
      NOR2_X1 XNOR_1_2_BUFF1_NUM188 (.ZN (N959), .A1 (XNOR_1_1_BUFF1_NUM188_OUT), .A2 (GND));
      wire XNOR_1_1_BUFF1_NUM189_OUT;
      NOR2_X1 XNOR_1_1_BUFF1_NUM189 (.ZN (XNOR_1_1_BUFF1_NUM189_OUT), .A1 (N574), .A2 (GND));
      NOR2_X1 XNOR_1_2_BUFF1_NUM189 (.ZN (N962), .A1 (XNOR_1_1_BUFF1_NUM189_OUT), .A2 (GND));
      wire XNOR_1_1_BUFF1_NUM190_OUT;
      NOR2_X1 XNOR_1_1_BUFF1_NUM190 (.ZN (XNOR_1_1_BUFF1_NUM190_OUT), .A1 (N580), .A2 (GND));
      NOR2_X1 XNOR_1_2_BUFF1_NUM190 (.ZN (N965), .A1 (XNOR_1_1_BUFF1_NUM190_OUT), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM191 (.ZN (N968), .A1 (N706), .A2 (GND));
      wire XNOR_1_1_BUFF1_NUM192_OUT;
      NOR2_X1 XNOR_1_1_BUFF1_NUM192 (.ZN (XNOR_1_1_BUFF1_NUM192_OUT), .A1 (N580), .A2 (GND));
      NOR2_X1 XNOR_1_2_BUFF1_NUM192 (.ZN (N969), .A1 (XNOR_1_1_BUFF1_NUM192_OUT), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM193 (.ZN (N972), .A1 (N709), .A2 (GND));
      wire XNOR_1_1_BUFF1_NUM194_OUT;
      NOR2_X1 XNOR_1_1_BUFF1_NUM194 (.ZN (XNOR_1_1_BUFF1_NUM194_OUT), .A1 (N586), .A2 (GND));
      NOR2_X1 XNOR_1_2_BUFF1_NUM194 (.ZN (N973), .A1 (XNOR_1_1_BUFF1_NUM194_OUT), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM195 (.ZN (N976), .A1 (N712), .A2 (GND));
      wire XNOR_1_1_BUFF1_NUM196_OUT;
      NOR2_X1 XNOR_1_1_BUFF1_NUM196 (.ZN (XNOR_1_1_BUFF1_NUM196_OUT), .A1 (N586), .A2 (GND));
      NOR2_X1 XNOR_1_2_BUFF1_NUM196 (.ZN (N977), .A1 (XNOR_1_1_BUFF1_NUM196_OUT), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM197 (.ZN (N980), .A1 (N715), .A2 (GND));
      wire XNOR_1_1_BUFF1_NUM198_OUT;
      NOR2_X1 XNOR_1_1_BUFF1_NUM198 (.ZN (XNOR_1_1_BUFF1_NUM198_OUT), .A1 (N592), .A2 (GND));
      NOR2_X1 XNOR_1_2_BUFF1_NUM198 (.ZN (N981), .A1 (XNOR_1_1_BUFF1_NUM198_OUT), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM199 (.ZN (N984), .A1 (N628), .A2 (GND));
      wire XNOR_1_1_BUFF1_NUM200_OUT;
      NOR2_X1 XNOR_1_1_BUFF1_NUM200 (.ZN (XNOR_1_1_BUFF1_NUM200_OUT), .A1 (N592), .A2 (GND));
      NOR2_X1 XNOR_1_2_BUFF1_NUM200 (.ZN (N985), .A1 (XNOR_1_1_BUFF1_NUM200_OUT), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM201 (.ZN (N988), .A1 (N718), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM202 (.ZN (N989), .A1 (N721), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM203 (.ZN (N990), .A1 (N634), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM204 (.ZN (N991), .A1 (N724), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM205 (.ZN (N992), .A1 (N727), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM206 (.ZN (N993), .A1 (N637), .A2 (GND));
      wire XNOR_1_1_BUFF1_NUM207_OUT;
      NOR2_X1 XNOR_1_1_BUFF1_NUM207 (.ZN (XNOR_1_1_BUFF1_NUM207_OUT), .A1 (N595), .A2 (GND));
      NOR2_X1 XNOR_1_2_BUFF1_NUM207 (.ZN (N994), .A1 (XNOR_1_1_BUFF1_NUM207_OUT), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM208 (.ZN (N997), .A1 (N730), .A2 (GND));
      wire XNOR_1_1_BUFF1_NUM209_OUT;
      NOR2_X1 XNOR_1_1_BUFF1_NUM209 (.ZN (XNOR_1_1_BUFF1_NUM209_OUT), .A1 (N595), .A2 (GND));
      NOR2_X1 XNOR_1_2_BUFF1_NUM209 (.ZN (N998), .A1 (XNOR_1_1_BUFF1_NUM209_OUT), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM210 (.ZN (N1001), .A1 (N733), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM211 (.ZN (N1002), .A1 (N736), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM212 (.ZN (N1003), .A1 (N739), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM213 (.ZN (N1004), .A1 (N640), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM214 (.ZN (N1005), .A1 (N742), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM215 (.ZN (N1006), .A1 (N745), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM216 (.ZN (N1007), .A1 (N646), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM217 (.ZN (N1008), .A1 (N748), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM218 (.ZN (N1009), .A1 (N751), .A2 (GND));
      wire XNOR_1_1_BUFF1_NUM219_OUT;
      NOR2_X1 XNOR_1_1_BUFF1_NUM219 (.ZN (XNOR_1_1_BUFF1_NUM219_OUT), .A1 (N559), .A2 (GND));
      NOR2_X1 XNOR_1_2_BUFF1_NUM219 (.ZN (N1010), .A1 (XNOR_1_1_BUFF1_NUM219_OUT), .A2 (GND));
      wire XNOR_1_1_BUFF1_NUM220_OUT;
      NOR2_X1 XNOR_1_1_BUFF1_NUM220 (.ZN (XNOR_1_1_BUFF1_NUM220_OUT), .A1 (N559), .A2 (GND));
      NOR2_X1 XNOR_1_2_BUFF1_NUM220 (.ZN (N1013), .A1 (XNOR_1_1_BUFF1_NUM220_OUT), .A2 (GND));
      wire XNOR_1_1_BUFF1_NUM221_OUT;
      NOR2_X1 XNOR_1_1_BUFF1_NUM221 (.ZN (XNOR_1_1_BUFF1_NUM221_OUT), .A1 (N565), .A2 (GND));
      NOR2_X1 XNOR_1_2_BUFF1_NUM221 (.ZN (N1016), .A1 (XNOR_1_1_BUFF1_NUM221_OUT), .A2 (GND));
      wire XNOR_1_1_BUFF1_NUM222_OUT;
      NOR2_X1 XNOR_1_1_BUFF1_NUM222 (.ZN (XNOR_1_1_BUFF1_NUM222_OUT), .A1 (N565), .A2 (GND));
      NOR2_X1 XNOR_1_2_BUFF1_NUM222 (.ZN (N1019), .A1 (XNOR_1_1_BUFF1_NUM222_OUT), .A2 (GND));
      wire XNOR_1_1_BUFF1_NUM223_OUT;
      NOR2_X1 XNOR_1_1_BUFF1_NUM223 (.ZN (XNOR_1_1_BUFF1_NUM223_OUT), .A1 (N571), .A2 (GND));
      NOR2_X1 XNOR_1_2_BUFF1_NUM223 (.ZN (N1022), .A1 (XNOR_1_1_BUFF1_NUM223_OUT), .A2 (GND));
      wire XNOR_1_1_BUFF1_NUM224_OUT;
      NOR2_X1 XNOR_1_1_BUFF1_NUM224 (.ZN (XNOR_1_1_BUFF1_NUM224_OUT), .A1 (N571), .A2 (GND));
      NOR2_X1 XNOR_1_2_BUFF1_NUM224 (.ZN (N1025), .A1 (XNOR_1_1_BUFF1_NUM224_OUT), .A2 (GND));
      wire XNOR_1_1_BUFF1_NUM225_OUT;
      NOR2_X1 XNOR_1_1_BUFF1_NUM225 (.ZN (XNOR_1_1_BUFF1_NUM225_OUT), .A1 (N577), .A2 (GND));
      NOR2_X1 XNOR_1_2_BUFF1_NUM225 (.ZN (N1028), .A1 (XNOR_1_1_BUFF1_NUM225_OUT), .A2 (GND));
      wire XNOR_1_1_BUFF1_NUM226_OUT;
      NOR2_X1 XNOR_1_1_BUFF1_NUM226 (.ZN (XNOR_1_1_BUFF1_NUM226_OUT), .A1 (N577), .A2 (GND));
      NOR2_X1 XNOR_1_2_BUFF1_NUM226 (.ZN (N1031), .A1 (XNOR_1_1_BUFF1_NUM226_OUT), .A2 (GND));
      wire XNOR_1_1_BUFF1_NUM227_OUT;
      NOR2_X1 XNOR_1_1_BUFF1_NUM227 (.ZN (XNOR_1_1_BUFF1_NUM227_OUT), .A1 (N583), .A2 (GND));
      NOR2_X1 XNOR_1_2_BUFF1_NUM227 (.ZN (N1034), .A1 (XNOR_1_1_BUFF1_NUM227_OUT), .A2 (GND));
      wire XNOR_1_1_BUFF1_NUM228_OUT;
      NOR2_X1 XNOR_1_1_BUFF1_NUM228 (.ZN (XNOR_1_1_BUFF1_NUM228_OUT), .A1 (N583), .A2 (GND));
      NOR2_X1 XNOR_1_2_BUFF1_NUM228 (.ZN (N1037), .A1 (XNOR_1_1_BUFF1_NUM228_OUT), .A2 (GND));
      wire XNOR_1_1_BUFF1_NUM229_OUT;
      NOR2_X1 XNOR_1_1_BUFF1_NUM229 (.ZN (XNOR_1_1_BUFF1_NUM229_OUT), .A1 (N589), .A2 (GND));
      NOR2_X1 XNOR_1_2_BUFF1_NUM229 (.ZN (N1040), .A1 (XNOR_1_1_BUFF1_NUM229_OUT), .A2 (GND));
      wire XNOR_1_1_BUFF1_NUM230_OUT;
      NOR2_X1 XNOR_1_1_BUFF1_NUM230 (.ZN (XNOR_1_1_BUFF1_NUM230_OUT), .A1 (N589), .A2 (GND));
      NOR2_X1 XNOR_1_2_BUFF1_NUM230 (.ZN (N1043), .A1 (XNOR_1_1_BUFF1_NUM230_OUT), .A2 (GND));
      wire XNOR_1_1_BUFF1_NUM231_OUT;
      NOR2_X1 XNOR_1_1_BUFF1_NUM231 (.ZN (XNOR_1_1_BUFF1_NUM231_OUT), .A1 (N598), .A2 (GND));
      NOR2_X1 XNOR_1_2_BUFF1_NUM231 (.ZN (N1046), .A1 (XNOR_1_1_BUFF1_NUM231_OUT), .A2 (GND));
      wire XNOR_1_1_BUFF1_NUM232_OUT;
      NOR2_X1 XNOR_1_1_BUFF1_NUM232 (.ZN (XNOR_1_1_BUFF1_NUM232_OUT), .A1 (N598), .A2 (GND));
      NOR2_X1 XNOR_1_2_BUFF1_NUM232 (.ZN (N1049), .A1 (XNOR_1_1_BUFF1_NUM232_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM233_OUT, XNOR_1_2_NAND2_NUM233_OUT, XNOR_1_3_NAND2_NUM233_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM233 (.ZN (XNOR_1_1_NAND2_NUM233_OUT), .A1 (N619), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM233 (.ZN (XNOR_1_2_NAND2_NUM233_OUT), .A1 (GND), .A2 (N888));
      NOR2_X1 XNOR_1_3_NAND2_NUM233 (.ZN (XNOR_1_3_NAND2_NUM233_OUT), .A1 (XNOR_1_1_NAND2_NUM233_OUT), .A2 (XNOR_1_2_NAND2_NUM233_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM233 (.ZN (N1054), .A1 (XNOR_1_3_NAND2_NUM233_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM234_OUT, XNOR_1_2_NAND2_NUM234_OUT, XNOR_1_3_NAND2_NUM234_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM234 (.ZN (XNOR_1_1_NAND2_NUM234_OUT), .A1 (N616), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM234 (.ZN (XNOR_1_2_NAND2_NUM234_OUT), .A1 (GND), .A2 (N889));
      NOR2_X1 XNOR_1_3_NAND2_NUM234 (.ZN (XNOR_1_3_NAND2_NUM234_OUT), .A1 (XNOR_1_1_NAND2_NUM234_OUT), .A2 (XNOR_1_2_NAND2_NUM234_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM234 (.ZN (N1055), .A1 (XNOR_1_3_NAND2_NUM234_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM235_OUT, XNOR_1_2_NAND2_NUM235_OUT, XNOR_1_3_NAND2_NUM235_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM235 (.ZN (XNOR_1_1_NAND2_NUM235_OUT), .A1 (N625), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM235 (.ZN (XNOR_1_2_NAND2_NUM235_OUT), .A1 (GND), .A2 (N890));
      NOR2_X1 XNOR_1_3_NAND2_NUM235 (.ZN (XNOR_1_3_NAND2_NUM235_OUT), .A1 (XNOR_1_1_NAND2_NUM235_OUT), .A2 (XNOR_1_2_NAND2_NUM235_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM235 (.ZN (N1063), .A1 (XNOR_1_3_NAND2_NUM235_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM236_OUT, XNOR_1_2_NAND2_NUM236_OUT, XNOR_1_3_NAND2_NUM236_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM236 (.ZN (XNOR_1_1_NAND2_NUM236_OUT), .A1 (N622), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM236 (.ZN (XNOR_1_2_NAND2_NUM236_OUT), .A1 (GND), .A2 (N891));
      NOR2_X1 XNOR_1_3_NAND2_NUM236 (.ZN (XNOR_1_3_NAND2_NUM236_OUT), .A1 (XNOR_1_1_NAND2_NUM236_OUT), .A2 (XNOR_1_2_NAND2_NUM236_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM236 (.ZN (N1064), .A1 (XNOR_1_3_NAND2_NUM236_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM237_OUT, XNOR_1_2_NAND2_NUM237_OUT, XNOR_1_3_NAND2_NUM237_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM237 (.ZN (XNOR_1_1_NAND2_NUM237_OUT), .A1 (N655), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM237 (.ZN (XNOR_1_2_NAND2_NUM237_OUT), .A1 (GND), .A2 (N895));
      NOR2_X1 XNOR_1_3_NAND2_NUM237 (.ZN (XNOR_1_3_NAND2_NUM237_OUT), .A1 (XNOR_1_1_NAND2_NUM237_OUT), .A2 (XNOR_1_2_NAND2_NUM237_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM237 (.ZN (N1067), .A1 (XNOR_1_3_NAND2_NUM237_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM238_OUT, XNOR_1_2_NAND2_NUM238_OUT, XNOR_1_3_NAND2_NUM238_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM238 (.ZN (XNOR_1_1_NAND2_NUM238_OUT), .A1 (N652), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM238 (.ZN (XNOR_1_2_NAND2_NUM238_OUT), .A1 (GND), .A2 (N896));
      NOR2_X1 XNOR_1_3_NAND2_NUM238 (.ZN (XNOR_1_3_NAND2_NUM238_OUT), .A1 (XNOR_1_1_NAND2_NUM238_OUT), .A2 (XNOR_1_2_NAND2_NUM238_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM238 (.ZN (N1068), .A1 (XNOR_1_3_NAND2_NUM238_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM239_OUT, XNOR_1_2_NAND2_NUM239_OUT, XNOR_1_3_NAND2_NUM239_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM239 (.ZN (XNOR_1_1_NAND2_NUM239_OUT), .A1 (N721), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM239 (.ZN (XNOR_1_2_NAND2_NUM239_OUT), .A1 (GND), .A2 (N988));
      NOR2_X1 XNOR_1_3_NAND2_NUM239 (.ZN (XNOR_1_3_NAND2_NUM239_OUT), .A1 (XNOR_1_1_NAND2_NUM239_OUT), .A2 (XNOR_1_2_NAND2_NUM239_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM239 (.ZN (N1119), .A1 (XNOR_1_3_NAND2_NUM239_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM240_OUT, XNOR_1_2_NAND2_NUM240_OUT, XNOR_1_3_NAND2_NUM240_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM240 (.ZN (XNOR_1_1_NAND2_NUM240_OUT), .A1 (N718), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM240 (.ZN (XNOR_1_2_NAND2_NUM240_OUT), .A1 (GND), .A2 (N989));
      NOR2_X1 XNOR_1_3_NAND2_NUM240 (.ZN (XNOR_1_3_NAND2_NUM240_OUT), .A1 (XNOR_1_1_NAND2_NUM240_OUT), .A2 (XNOR_1_2_NAND2_NUM240_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM240 (.ZN (N1120), .A1 (XNOR_1_3_NAND2_NUM240_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM241_OUT, XNOR_1_2_NAND2_NUM241_OUT, XNOR_1_3_NAND2_NUM241_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM241 (.ZN (XNOR_1_1_NAND2_NUM241_OUT), .A1 (N727), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM241 (.ZN (XNOR_1_2_NAND2_NUM241_OUT), .A1 (GND), .A2 (N991));
      NOR2_X1 XNOR_1_3_NAND2_NUM241 (.ZN (XNOR_1_3_NAND2_NUM241_OUT), .A1 (XNOR_1_1_NAND2_NUM241_OUT), .A2 (XNOR_1_2_NAND2_NUM241_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM241 (.ZN (N1121), .A1 (XNOR_1_3_NAND2_NUM241_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM242_OUT, XNOR_1_2_NAND2_NUM242_OUT, XNOR_1_3_NAND2_NUM242_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM242 (.ZN (XNOR_1_1_NAND2_NUM242_OUT), .A1 (N724), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM242 (.ZN (XNOR_1_2_NAND2_NUM242_OUT), .A1 (GND), .A2 (N992));
      NOR2_X1 XNOR_1_3_NAND2_NUM242 (.ZN (XNOR_1_3_NAND2_NUM242_OUT), .A1 (XNOR_1_1_NAND2_NUM242_OUT), .A2 (XNOR_1_2_NAND2_NUM242_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM242 (.ZN (N1122), .A1 (XNOR_1_3_NAND2_NUM242_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM243_OUT, XNOR_1_2_NAND2_NUM243_OUT, XNOR_1_3_NAND2_NUM243_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM243 (.ZN (XNOR_1_1_NAND2_NUM243_OUT), .A1 (N739), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM243 (.ZN (XNOR_1_2_NAND2_NUM243_OUT), .A1 (GND), .A2 (N1002));
      NOR2_X1 XNOR_1_3_NAND2_NUM243 (.ZN (XNOR_1_3_NAND2_NUM243_OUT), .A1 (XNOR_1_1_NAND2_NUM243_OUT), .A2 (XNOR_1_2_NAND2_NUM243_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM243 (.ZN (N1128), .A1 (XNOR_1_3_NAND2_NUM243_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM244_OUT, XNOR_1_2_NAND2_NUM244_OUT, XNOR_1_3_NAND2_NUM244_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM244 (.ZN (XNOR_1_1_NAND2_NUM244_OUT), .A1 (N736), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM244 (.ZN (XNOR_1_2_NAND2_NUM244_OUT), .A1 (GND), .A2 (N1003));
      NOR2_X1 XNOR_1_3_NAND2_NUM244 (.ZN (XNOR_1_3_NAND2_NUM244_OUT), .A1 (XNOR_1_1_NAND2_NUM244_OUT), .A2 (XNOR_1_2_NAND2_NUM244_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM244 (.ZN (N1129), .A1 (XNOR_1_3_NAND2_NUM244_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM245_OUT, XNOR_1_2_NAND2_NUM245_OUT, XNOR_1_3_NAND2_NUM245_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM245 (.ZN (XNOR_1_1_NAND2_NUM245_OUT), .A1 (N745), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM245 (.ZN (XNOR_1_2_NAND2_NUM245_OUT), .A1 (GND), .A2 (N1005));
      NOR2_X1 XNOR_1_3_NAND2_NUM245 (.ZN (XNOR_1_3_NAND2_NUM245_OUT), .A1 (XNOR_1_1_NAND2_NUM245_OUT), .A2 (XNOR_1_2_NAND2_NUM245_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM245 (.ZN (N1130), .A1 (XNOR_1_3_NAND2_NUM245_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM246_OUT, XNOR_1_2_NAND2_NUM246_OUT, XNOR_1_3_NAND2_NUM246_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM246 (.ZN (XNOR_1_1_NAND2_NUM246_OUT), .A1 (N742), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM246 (.ZN (XNOR_1_2_NAND2_NUM246_OUT), .A1 (GND), .A2 (N1006));
      NOR2_X1 XNOR_1_3_NAND2_NUM246 (.ZN (XNOR_1_3_NAND2_NUM246_OUT), .A1 (XNOR_1_1_NAND2_NUM246_OUT), .A2 (XNOR_1_2_NAND2_NUM246_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM246 (.ZN (N1131), .A1 (XNOR_1_3_NAND2_NUM246_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM247_OUT, XNOR_1_2_NAND2_NUM247_OUT, XNOR_1_3_NAND2_NUM247_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM247 (.ZN (XNOR_1_1_NAND2_NUM247_OUT), .A1 (N751), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM247 (.ZN (XNOR_1_2_NAND2_NUM247_OUT), .A1 (GND), .A2 (N1008));
      NOR2_X1 XNOR_1_3_NAND2_NUM247 (.ZN (XNOR_1_3_NAND2_NUM247_OUT), .A1 (XNOR_1_1_NAND2_NUM247_OUT), .A2 (XNOR_1_2_NAND2_NUM247_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM247 (.ZN (N1132), .A1 (XNOR_1_3_NAND2_NUM247_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM248_OUT, XNOR_1_2_NAND2_NUM248_OUT, XNOR_1_3_NAND2_NUM248_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM248 (.ZN (XNOR_1_1_NAND2_NUM248_OUT), .A1 (N748), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM248 (.ZN (XNOR_1_2_NAND2_NUM248_OUT), .A1 (GND), .A2 (N1009));
      NOR2_X1 XNOR_1_3_NAND2_NUM248 (.ZN (XNOR_1_3_NAND2_NUM248_OUT), .A1 (XNOR_1_1_NAND2_NUM248_OUT), .A2 (XNOR_1_2_NAND2_NUM248_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM248 (.ZN (N1133), .A1 (XNOR_1_3_NAND2_NUM248_OUT), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM249 (.ZN (N1148), .A1 (N939), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM250 (.ZN (N1149), .A1 (N935), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM251_OUT, XNOR_1_2_NAND2_NUM251_OUT, XNOR_1_3_NAND2_NUM251_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM251 (.ZN (XNOR_1_1_NAND2_NUM251_OUT), .A1 (N1054), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM251 (.ZN (XNOR_1_2_NAND2_NUM251_OUT), .A1 (GND), .A2 (N1055));
      NOR2_X1 XNOR_1_3_NAND2_NUM251 (.ZN (XNOR_1_3_NAND2_NUM251_OUT), .A1 (XNOR_1_1_NAND2_NUM251_OUT), .A2 (XNOR_1_2_NAND2_NUM251_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM251 (.ZN (N1150), .A1 (XNOR_1_3_NAND2_NUM251_OUT), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM252 (.ZN (N1151), .A1 (N943), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM253 (.ZN (N1152), .A1 (N947), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM254 (.ZN (N1153), .A1 (N955), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM255 (.ZN (N1154), .A1 (N951), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM256 (.ZN (N1155), .A1 (N962), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM257 (.ZN (N1156), .A1 (N969), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM258 (.ZN (N1157), .A1 (N977), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM259_OUT, XNOR_1_2_NAND2_NUM259_OUT, XNOR_1_3_NAND2_NUM259_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM259 (.ZN (XNOR_1_1_NAND2_NUM259_OUT), .A1 (N1063), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM259 (.ZN (XNOR_1_2_NAND2_NUM259_OUT), .A1 (GND), .A2 (N1064));
      NOR2_X1 XNOR_1_3_NAND2_NUM259 (.ZN (XNOR_1_3_NAND2_NUM259_OUT), .A1 (XNOR_1_1_NAND2_NUM259_OUT), .A2 (XNOR_1_2_NAND2_NUM259_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM259 (.ZN (N1158), .A1 (XNOR_1_3_NAND2_NUM259_OUT), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM260 (.ZN (N1159), .A1 (N985), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM261_OUT, XNOR_1_2_NAND2_NUM261_OUT, XNOR_1_3_NAND2_NUM261_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM261 (.ZN (XNOR_1_1_NAND2_NUM261_OUT), .A1 (N985), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM261 (.ZN (XNOR_1_2_NAND2_NUM261_OUT), .A1 (GND), .A2 (N892));
      NOR2_X1 XNOR_1_3_NAND2_NUM261 (.ZN (XNOR_1_3_NAND2_NUM261_OUT), .A1 (XNOR_1_1_NAND2_NUM261_OUT), .A2 (XNOR_1_2_NAND2_NUM261_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM261 (.ZN (N1160), .A1 (XNOR_1_3_NAND2_NUM261_OUT), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM262 (.ZN (N1161), .A1 (N998), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM263_OUT, XNOR_1_2_NAND2_NUM263_OUT, XNOR_1_3_NAND2_NUM263_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM263 (.ZN (XNOR_1_1_NAND2_NUM263_OUT), .A1 (N1067), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM263 (.ZN (XNOR_1_2_NAND2_NUM263_OUT), .A1 (GND), .A2 (N1068));
      NOR2_X1 XNOR_1_3_NAND2_NUM263 (.ZN (XNOR_1_3_NAND2_NUM263_OUT), .A1 (XNOR_1_1_NAND2_NUM263_OUT), .A2 (XNOR_1_2_NAND2_NUM263_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM263 (.ZN (N1162), .A1 (XNOR_1_3_NAND2_NUM263_OUT), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM264 (.ZN (N1163), .A1 (N899), .A2 (GND));
      wire XNOR_1_1_BUFF1_NUM265_OUT;
      NOR2_X1 XNOR_1_1_BUFF1_NUM265 (.ZN (XNOR_1_1_BUFF1_NUM265_OUT), .A1 (N899), .A2 (GND));
      NOR2_X1 XNOR_1_2_BUFF1_NUM265 (.ZN (N1164), .A1 (XNOR_1_1_BUFF1_NUM265_OUT), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM266 (.ZN (N1167), .A1 (N903), .A2 (GND));
      wire XNOR_1_1_BUFF1_NUM267_OUT;
      NOR2_X1 XNOR_1_1_BUFF1_NUM267 (.ZN (XNOR_1_1_BUFF1_NUM267_OUT), .A1 (N903), .A2 (GND));
      NOR2_X1 XNOR_1_2_BUFF1_NUM267 (.ZN (N1168), .A1 (XNOR_1_1_BUFF1_NUM267_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM268_OUT, XNOR_1_2_NAND2_NUM268_OUT, XNOR_1_3_NAND2_NUM268_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM268 (.ZN (XNOR_1_1_NAND2_NUM268_OUT), .A1 (N921), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM268 (.ZN (XNOR_1_2_NAND2_NUM268_OUT), .A1 (GND), .A2 (N923));
      NOR2_X1 XNOR_1_3_NAND2_NUM268 (.ZN (XNOR_1_3_NAND2_NUM268_OUT), .A1 (XNOR_1_1_NAND2_NUM268_OUT), .A2 (XNOR_1_2_NAND2_NUM268_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM268 (.ZN (N1171), .A1 (XNOR_1_3_NAND2_NUM268_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM269_OUT, XNOR_1_2_NAND2_NUM269_OUT, XNOR_1_3_NAND2_NUM269_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM269 (.ZN (XNOR_1_1_NAND2_NUM269_OUT), .A1 (N922), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM269 (.ZN (XNOR_1_2_NAND2_NUM269_OUT), .A1 (GND), .A2 (N923));
      NOR2_X1 XNOR_1_3_NAND2_NUM269 (.ZN (XNOR_1_3_NAND2_NUM269_OUT), .A1 (XNOR_1_1_NAND2_NUM269_OUT), .A2 (XNOR_1_2_NAND2_NUM269_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM269 (.ZN (N1188), .A1 (XNOR_1_3_NAND2_NUM269_OUT), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM270 (.ZN (N1205), .A1 (N1010), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM271_OUT, XNOR_1_2_NAND2_NUM271_OUT, XNOR_1_3_NAND2_NUM271_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM271 (.ZN (XNOR_1_1_NAND2_NUM271_OUT), .A1 (N1010), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM271 (.ZN (XNOR_1_2_NAND2_NUM271_OUT), .A1 (GND), .A2 (N938));
      NOR2_X1 XNOR_1_3_NAND2_NUM271 (.ZN (XNOR_1_3_NAND2_NUM271_OUT), .A1 (XNOR_1_1_NAND2_NUM271_OUT), .A2 (XNOR_1_2_NAND2_NUM271_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM271 (.ZN (N1206), .A1 (XNOR_1_3_NAND2_NUM271_OUT), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM272 (.ZN (N1207), .A1 (N1013), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM273_OUT, XNOR_1_2_NAND2_NUM273_OUT, XNOR_1_3_NAND2_NUM273_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM273 (.ZN (XNOR_1_1_NAND2_NUM273_OUT), .A1 (N1013), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM273 (.ZN (XNOR_1_2_NAND2_NUM273_OUT), .A1 (GND), .A2 (N942));
      NOR2_X1 XNOR_1_3_NAND2_NUM273 (.ZN (XNOR_1_3_NAND2_NUM273_OUT), .A1 (XNOR_1_1_NAND2_NUM273_OUT), .A2 (XNOR_1_2_NAND2_NUM273_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM273 (.ZN (N1208), .A1 (XNOR_1_3_NAND2_NUM273_OUT), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM274 (.ZN (N1209), .A1 (N1016), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM275_OUT, XNOR_1_2_NAND2_NUM275_OUT, XNOR_1_3_NAND2_NUM275_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM275 (.ZN (XNOR_1_1_NAND2_NUM275_OUT), .A1 (N1016), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM275 (.ZN (XNOR_1_2_NAND2_NUM275_OUT), .A1 (GND), .A2 (N946));
      NOR2_X1 XNOR_1_3_NAND2_NUM275 (.ZN (XNOR_1_3_NAND2_NUM275_OUT), .A1 (XNOR_1_1_NAND2_NUM275_OUT), .A2 (XNOR_1_2_NAND2_NUM275_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM275 (.ZN (N1210), .A1 (XNOR_1_3_NAND2_NUM275_OUT), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM276 (.ZN (N1211), .A1 (N1019), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM277_OUT, XNOR_1_2_NAND2_NUM277_OUT, XNOR_1_3_NAND2_NUM277_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM277 (.ZN (XNOR_1_1_NAND2_NUM277_OUT), .A1 (N1019), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM277 (.ZN (XNOR_1_2_NAND2_NUM277_OUT), .A1 (GND), .A2 (N950));
      NOR2_X1 XNOR_1_3_NAND2_NUM277 (.ZN (XNOR_1_3_NAND2_NUM277_OUT), .A1 (XNOR_1_1_NAND2_NUM277_OUT), .A2 (XNOR_1_2_NAND2_NUM277_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM277 (.ZN (N1212), .A1 (XNOR_1_3_NAND2_NUM277_OUT), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM278 (.ZN (N1213), .A1 (N1022), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM279_OUT, XNOR_1_2_NAND2_NUM279_OUT, XNOR_1_3_NAND2_NUM279_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM279 (.ZN (XNOR_1_1_NAND2_NUM279_OUT), .A1 (N1022), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM279 (.ZN (XNOR_1_2_NAND2_NUM279_OUT), .A1 (GND), .A2 (N954));
      NOR2_X1 XNOR_1_3_NAND2_NUM279 (.ZN (XNOR_1_3_NAND2_NUM279_OUT), .A1 (XNOR_1_1_NAND2_NUM279_OUT), .A2 (XNOR_1_2_NAND2_NUM279_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM279 (.ZN (N1214), .A1 (XNOR_1_3_NAND2_NUM279_OUT), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM280 (.ZN (N1215), .A1 (N1025), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM281_OUT, XNOR_1_2_NAND2_NUM281_OUT, XNOR_1_3_NAND2_NUM281_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM281 (.ZN (XNOR_1_1_NAND2_NUM281_OUT), .A1 (N1025), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM281 (.ZN (XNOR_1_2_NAND2_NUM281_OUT), .A1 (GND), .A2 (N958));
      NOR2_X1 XNOR_1_3_NAND2_NUM281 (.ZN (XNOR_1_3_NAND2_NUM281_OUT), .A1 (XNOR_1_1_NAND2_NUM281_OUT), .A2 (XNOR_1_2_NAND2_NUM281_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM281 (.ZN (N1216), .A1 (XNOR_1_3_NAND2_NUM281_OUT), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM282 (.ZN (N1217), .A1 (N1028), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM283 (.ZN (N1218), .A1 (N959), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM284 (.ZN (N1219), .A1 (N1031), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM285 (.ZN (N1220), .A1 (N1034), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM286_OUT, XNOR_1_2_NAND2_NUM286_OUT, XNOR_1_3_NAND2_NUM286_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM286 (.ZN (XNOR_1_1_NAND2_NUM286_OUT), .A1 (N1034), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM286 (.ZN (XNOR_1_2_NAND2_NUM286_OUT), .A1 (GND), .A2 (N968));
      NOR2_X1 XNOR_1_3_NAND2_NUM286 (.ZN (XNOR_1_3_NAND2_NUM286_OUT), .A1 (XNOR_1_1_NAND2_NUM286_OUT), .A2 (XNOR_1_2_NAND2_NUM286_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM286 (.ZN (N1221), .A1 (XNOR_1_3_NAND2_NUM286_OUT), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM287 (.ZN (N1222), .A1 (N965), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM288 (.ZN (N1223), .A1 (N1037), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM289_OUT, XNOR_1_2_NAND2_NUM289_OUT, XNOR_1_3_NAND2_NUM289_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM289 (.ZN (XNOR_1_1_NAND2_NUM289_OUT), .A1 (N1037), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM289 (.ZN (XNOR_1_2_NAND2_NUM289_OUT), .A1 (GND), .A2 (N972));
      NOR2_X1 XNOR_1_3_NAND2_NUM289 (.ZN (XNOR_1_3_NAND2_NUM289_OUT), .A1 (XNOR_1_1_NAND2_NUM289_OUT), .A2 (XNOR_1_2_NAND2_NUM289_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM289 (.ZN (N1224), .A1 (XNOR_1_3_NAND2_NUM289_OUT), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM290 (.ZN (N1225), .A1 (N1040), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM291_OUT, XNOR_1_2_NAND2_NUM291_OUT, XNOR_1_3_NAND2_NUM291_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM291 (.ZN (XNOR_1_1_NAND2_NUM291_OUT), .A1 (N1040), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM291 (.ZN (XNOR_1_2_NAND2_NUM291_OUT), .A1 (GND), .A2 (N976));
      NOR2_X1 XNOR_1_3_NAND2_NUM291 (.ZN (XNOR_1_3_NAND2_NUM291_OUT), .A1 (XNOR_1_1_NAND2_NUM291_OUT), .A2 (XNOR_1_2_NAND2_NUM291_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM291 (.ZN (N1226), .A1 (XNOR_1_3_NAND2_NUM291_OUT), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM292 (.ZN (N1227), .A1 (N973), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM293 (.ZN (N1228), .A1 (N1043), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM294_OUT, XNOR_1_2_NAND2_NUM294_OUT, XNOR_1_3_NAND2_NUM294_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM294 (.ZN (XNOR_1_1_NAND2_NUM294_OUT), .A1 (N1043), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM294 (.ZN (XNOR_1_2_NAND2_NUM294_OUT), .A1 (GND), .A2 (N980));
      NOR2_X1 XNOR_1_3_NAND2_NUM294 (.ZN (XNOR_1_3_NAND2_NUM294_OUT), .A1 (XNOR_1_1_NAND2_NUM294_OUT), .A2 (XNOR_1_2_NAND2_NUM294_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM294 (.ZN (N1229), .A1 (XNOR_1_3_NAND2_NUM294_OUT), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM295 (.ZN (N1230), .A1 (N981), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM296_OUT, XNOR_1_2_NAND2_NUM296_OUT, XNOR_1_3_NAND2_NUM296_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM296 (.ZN (XNOR_1_1_NAND2_NUM296_OUT), .A1 (N981), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM296 (.ZN (XNOR_1_2_NAND2_NUM296_OUT), .A1 (GND), .A2 (N984));
      NOR2_X1 XNOR_1_3_NAND2_NUM296 (.ZN (XNOR_1_3_NAND2_NUM296_OUT), .A1 (XNOR_1_1_NAND2_NUM296_OUT), .A2 (XNOR_1_2_NAND2_NUM296_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM296 (.ZN (N1231), .A1 (XNOR_1_3_NAND2_NUM296_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM297_OUT, XNOR_1_2_NAND2_NUM297_OUT, XNOR_1_3_NAND2_NUM297_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM297 (.ZN (XNOR_1_1_NAND2_NUM297_OUT), .A1 (N1119), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM297 (.ZN (XNOR_1_2_NAND2_NUM297_OUT), .A1 (GND), .A2 (N1120));
      NOR2_X1 XNOR_1_3_NAND2_NUM297 (.ZN (XNOR_1_3_NAND2_NUM297_OUT), .A1 (XNOR_1_1_NAND2_NUM297_OUT), .A2 (XNOR_1_2_NAND2_NUM297_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM297 (.ZN (N1232), .A1 (XNOR_1_3_NAND2_NUM297_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM298_OUT, XNOR_1_2_NAND2_NUM298_OUT, XNOR_1_3_NAND2_NUM298_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM298 (.ZN (XNOR_1_1_NAND2_NUM298_OUT), .A1 (N1121), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM298 (.ZN (XNOR_1_2_NAND2_NUM298_OUT), .A1 (GND), .A2 (N1122));
      NOR2_X1 XNOR_1_3_NAND2_NUM298 (.ZN (XNOR_1_3_NAND2_NUM298_OUT), .A1 (XNOR_1_1_NAND2_NUM298_OUT), .A2 (XNOR_1_2_NAND2_NUM298_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM298 (.ZN (N1235), .A1 (XNOR_1_3_NAND2_NUM298_OUT), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM299 (.ZN (N1238), .A1 (N1046), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM300_OUT, XNOR_1_2_NAND2_NUM300_OUT, XNOR_1_3_NAND2_NUM300_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM300 (.ZN (XNOR_1_1_NAND2_NUM300_OUT), .A1 (N1046), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM300 (.ZN (XNOR_1_2_NAND2_NUM300_OUT), .A1 (GND), .A2 (N997));
      NOR2_X1 XNOR_1_3_NAND2_NUM300 (.ZN (XNOR_1_3_NAND2_NUM300_OUT), .A1 (XNOR_1_1_NAND2_NUM300_OUT), .A2 (XNOR_1_2_NAND2_NUM300_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM300 (.ZN (N1239), .A1 (XNOR_1_3_NAND2_NUM300_OUT), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM301 (.ZN (N1240), .A1 (N994), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM302 (.ZN (N1241), .A1 (N1049), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM303_OUT, XNOR_1_2_NAND2_NUM303_OUT, XNOR_1_3_NAND2_NUM303_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM303 (.ZN (XNOR_1_1_NAND2_NUM303_OUT), .A1 (N1049), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM303 (.ZN (XNOR_1_2_NAND2_NUM303_OUT), .A1 (GND), .A2 (N1001));
      NOR2_X1 XNOR_1_3_NAND2_NUM303 (.ZN (XNOR_1_3_NAND2_NUM303_OUT), .A1 (XNOR_1_1_NAND2_NUM303_OUT), .A2 (XNOR_1_2_NAND2_NUM303_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM303 (.ZN (N1242), .A1 (XNOR_1_3_NAND2_NUM303_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM304_OUT, XNOR_1_2_NAND2_NUM304_OUT, XNOR_1_3_NAND2_NUM304_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM304 (.ZN (XNOR_1_1_NAND2_NUM304_OUT), .A1 (N1128), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM304 (.ZN (XNOR_1_2_NAND2_NUM304_OUT), .A1 (GND), .A2 (N1129));
      NOR2_X1 XNOR_1_3_NAND2_NUM304 (.ZN (XNOR_1_3_NAND2_NUM304_OUT), .A1 (XNOR_1_1_NAND2_NUM304_OUT), .A2 (XNOR_1_2_NAND2_NUM304_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM304 (.ZN (N1243), .A1 (XNOR_1_3_NAND2_NUM304_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM305_OUT, XNOR_1_2_NAND2_NUM305_OUT, XNOR_1_3_NAND2_NUM305_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM305 (.ZN (XNOR_1_1_NAND2_NUM305_OUT), .A1 (N1130), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM305 (.ZN (XNOR_1_2_NAND2_NUM305_OUT), .A1 (GND), .A2 (N1131));
      NOR2_X1 XNOR_1_3_NAND2_NUM305 (.ZN (XNOR_1_3_NAND2_NUM305_OUT), .A1 (XNOR_1_1_NAND2_NUM305_OUT), .A2 (XNOR_1_2_NAND2_NUM305_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM305 (.ZN (N1246), .A1 (XNOR_1_3_NAND2_NUM305_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM306_OUT, XNOR_1_2_NAND2_NUM306_OUT, XNOR_1_3_NAND2_NUM306_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM306 (.ZN (XNOR_1_1_NAND2_NUM306_OUT), .A1 (N1132), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM306 (.ZN (XNOR_1_2_NAND2_NUM306_OUT), .A1 (GND), .A2 (N1133));
      NOR2_X1 XNOR_1_3_NAND2_NUM306 (.ZN (XNOR_1_3_NAND2_NUM306_OUT), .A1 (XNOR_1_1_NAND2_NUM306_OUT), .A2 (XNOR_1_2_NAND2_NUM306_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM306 (.ZN (N1249), .A1 (XNOR_1_3_NAND2_NUM306_OUT), .A2 (GND));
      wire XNOR_1_1_BUFF1_NUM307_OUT;
      NOR2_X1 XNOR_1_1_BUFF1_NUM307 (.ZN (XNOR_1_1_BUFF1_NUM307_OUT), .A1 (N907), .A2 (GND));
      NOR2_X1 XNOR_1_2_BUFF1_NUM307 (.ZN (N1252), .A1 (XNOR_1_1_BUFF1_NUM307_OUT), .A2 (GND));
      wire XNOR_1_1_BUFF1_NUM308_OUT;
      NOR2_X1 XNOR_1_1_BUFF1_NUM308 (.ZN (XNOR_1_1_BUFF1_NUM308_OUT), .A1 (N907), .A2 (GND));
      NOR2_X1 XNOR_1_2_BUFF1_NUM308 (.ZN (N1255), .A1 (XNOR_1_1_BUFF1_NUM308_OUT), .A2 (GND));
      wire XNOR_1_1_BUFF1_NUM309_OUT;
      NOR2_X1 XNOR_1_1_BUFF1_NUM309 (.ZN (XNOR_1_1_BUFF1_NUM309_OUT), .A1 (N910), .A2 (GND));
      NOR2_X1 XNOR_1_2_BUFF1_NUM309 (.ZN (N1258), .A1 (XNOR_1_1_BUFF1_NUM309_OUT), .A2 (GND));
      wire XNOR_1_1_BUFF1_NUM310_OUT;
      NOR2_X1 XNOR_1_1_BUFF1_NUM310 (.ZN (XNOR_1_1_BUFF1_NUM310_OUT), .A1 (N910), .A2 (GND));
      NOR2_X1 XNOR_1_2_BUFF1_NUM310 (.ZN (N1261), .A1 (XNOR_1_1_BUFF1_NUM310_OUT), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM311 (.ZN (N1264), .A1 (N1150), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM312_OUT, XNOR_1_2_NAND2_NUM312_OUT, XNOR_1_3_NAND2_NUM312_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM312 (.ZN (XNOR_1_1_NAND2_NUM312_OUT), .A1 (N631), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM312 (.ZN (XNOR_1_2_NAND2_NUM312_OUT), .A1 (GND), .A2 (N1159));
      NOR2_X1 XNOR_1_3_NAND2_NUM312 (.ZN (XNOR_1_3_NAND2_NUM312_OUT), .A1 (XNOR_1_1_NAND2_NUM312_OUT), .A2 (XNOR_1_2_NAND2_NUM312_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM312 (.ZN (N1267), .A1 (XNOR_1_3_NAND2_NUM312_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM313_OUT, XNOR_1_2_NAND2_NUM313_OUT, XNOR_1_3_NAND2_NUM313_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM313 (.ZN (XNOR_1_1_NAND2_NUM313_OUT), .A1 (N688), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM313 (.ZN (XNOR_1_2_NAND2_NUM313_OUT), .A1 (GND), .A2 (N1205));
      NOR2_X1 XNOR_1_3_NAND2_NUM313 (.ZN (XNOR_1_3_NAND2_NUM313_OUT), .A1 (XNOR_1_1_NAND2_NUM313_OUT), .A2 (XNOR_1_2_NAND2_NUM313_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM313 (.ZN (N1309), .A1 (XNOR_1_3_NAND2_NUM313_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM314_OUT, XNOR_1_2_NAND2_NUM314_OUT, XNOR_1_3_NAND2_NUM314_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM314 (.ZN (XNOR_1_1_NAND2_NUM314_OUT), .A1 (N691), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM314 (.ZN (XNOR_1_2_NAND2_NUM314_OUT), .A1 (GND), .A2 (N1207));
      NOR2_X1 XNOR_1_3_NAND2_NUM314 (.ZN (XNOR_1_3_NAND2_NUM314_OUT), .A1 (XNOR_1_1_NAND2_NUM314_OUT), .A2 (XNOR_1_2_NAND2_NUM314_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM314 (.ZN (N1310), .A1 (XNOR_1_3_NAND2_NUM314_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM315_OUT, XNOR_1_2_NAND2_NUM315_OUT, XNOR_1_3_NAND2_NUM315_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM315 (.ZN (XNOR_1_1_NAND2_NUM315_OUT), .A1 (N694), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM315 (.ZN (XNOR_1_2_NAND2_NUM315_OUT), .A1 (GND), .A2 (N1209));
      NOR2_X1 XNOR_1_3_NAND2_NUM315 (.ZN (XNOR_1_3_NAND2_NUM315_OUT), .A1 (XNOR_1_1_NAND2_NUM315_OUT), .A2 (XNOR_1_2_NAND2_NUM315_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM315 (.ZN (N1311), .A1 (XNOR_1_3_NAND2_NUM315_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM316_OUT, XNOR_1_2_NAND2_NUM316_OUT, XNOR_1_3_NAND2_NUM316_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM316 (.ZN (XNOR_1_1_NAND2_NUM316_OUT), .A1 (N697), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM316 (.ZN (XNOR_1_2_NAND2_NUM316_OUT), .A1 (GND), .A2 (N1211));
      NOR2_X1 XNOR_1_3_NAND2_NUM316 (.ZN (XNOR_1_3_NAND2_NUM316_OUT), .A1 (XNOR_1_1_NAND2_NUM316_OUT), .A2 (XNOR_1_2_NAND2_NUM316_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM316 (.ZN (N1312), .A1 (XNOR_1_3_NAND2_NUM316_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM317_OUT, XNOR_1_2_NAND2_NUM317_OUT, XNOR_1_3_NAND2_NUM317_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM317 (.ZN (XNOR_1_1_NAND2_NUM317_OUT), .A1 (N700), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM317 (.ZN (XNOR_1_2_NAND2_NUM317_OUT), .A1 (GND), .A2 (N1213));
      NOR2_X1 XNOR_1_3_NAND2_NUM317 (.ZN (XNOR_1_3_NAND2_NUM317_OUT), .A1 (XNOR_1_1_NAND2_NUM317_OUT), .A2 (XNOR_1_2_NAND2_NUM317_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM317 (.ZN (N1313), .A1 (XNOR_1_3_NAND2_NUM317_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM318_OUT, XNOR_1_2_NAND2_NUM318_OUT, XNOR_1_3_NAND2_NUM318_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM318 (.ZN (XNOR_1_1_NAND2_NUM318_OUT), .A1 (N703), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM318 (.ZN (XNOR_1_2_NAND2_NUM318_OUT), .A1 (GND), .A2 (N1215));
      NOR2_X1 XNOR_1_3_NAND2_NUM318 (.ZN (XNOR_1_3_NAND2_NUM318_OUT), .A1 (XNOR_1_1_NAND2_NUM318_OUT), .A2 (XNOR_1_2_NAND2_NUM318_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM318 (.ZN (N1314), .A1 (XNOR_1_3_NAND2_NUM318_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM319_OUT, XNOR_1_2_NAND2_NUM319_OUT, XNOR_1_3_NAND2_NUM319_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM319 (.ZN (XNOR_1_1_NAND2_NUM319_OUT), .A1 (N706), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM319 (.ZN (XNOR_1_2_NAND2_NUM319_OUT), .A1 (GND), .A2 (N1220));
      NOR2_X1 XNOR_1_3_NAND2_NUM319 (.ZN (XNOR_1_3_NAND2_NUM319_OUT), .A1 (XNOR_1_1_NAND2_NUM319_OUT), .A2 (XNOR_1_2_NAND2_NUM319_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM319 (.ZN (N1315), .A1 (XNOR_1_3_NAND2_NUM319_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM320_OUT, XNOR_1_2_NAND2_NUM320_OUT, XNOR_1_3_NAND2_NUM320_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM320 (.ZN (XNOR_1_1_NAND2_NUM320_OUT), .A1 (N709), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM320 (.ZN (XNOR_1_2_NAND2_NUM320_OUT), .A1 (GND), .A2 (N1223));
      NOR2_X1 XNOR_1_3_NAND2_NUM320 (.ZN (XNOR_1_3_NAND2_NUM320_OUT), .A1 (XNOR_1_1_NAND2_NUM320_OUT), .A2 (XNOR_1_2_NAND2_NUM320_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM320 (.ZN (N1316), .A1 (XNOR_1_3_NAND2_NUM320_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM321_OUT, XNOR_1_2_NAND2_NUM321_OUT, XNOR_1_3_NAND2_NUM321_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM321 (.ZN (XNOR_1_1_NAND2_NUM321_OUT), .A1 (N712), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM321 (.ZN (XNOR_1_2_NAND2_NUM321_OUT), .A1 (GND), .A2 (N1225));
      NOR2_X1 XNOR_1_3_NAND2_NUM321 (.ZN (XNOR_1_3_NAND2_NUM321_OUT), .A1 (XNOR_1_1_NAND2_NUM321_OUT), .A2 (XNOR_1_2_NAND2_NUM321_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM321 (.ZN (N1317), .A1 (XNOR_1_3_NAND2_NUM321_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM322_OUT, XNOR_1_2_NAND2_NUM322_OUT, XNOR_1_3_NAND2_NUM322_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM322 (.ZN (XNOR_1_1_NAND2_NUM322_OUT), .A1 (N715), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM322 (.ZN (XNOR_1_2_NAND2_NUM322_OUT), .A1 (GND), .A2 (N1228));
      NOR2_X1 XNOR_1_3_NAND2_NUM322 (.ZN (XNOR_1_3_NAND2_NUM322_OUT), .A1 (XNOR_1_1_NAND2_NUM322_OUT), .A2 (XNOR_1_2_NAND2_NUM322_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM322 (.ZN (N1318), .A1 (XNOR_1_3_NAND2_NUM322_OUT), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM323 (.ZN (N1319), .A1 (N1158), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM324_OUT, XNOR_1_2_NAND2_NUM324_OUT, XNOR_1_3_NAND2_NUM324_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM324 (.ZN (XNOR_1_1_NAND2_NUM324_OUT), .A1 (N628), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM324 (.ZN (XNOR_1_2_NAND2_NUM324_OUT), .A1 (GND), .A2 (N1230));
      NOR2_X1 XNOR_1_3_NAND2_NUM324 (.ZN (XNOR_1_3_NAND2_NUM324_OUT), .A1 (XNOR_1_1_NAND2_NUM324_OUT), .A2 (XNOR_1_2_NAND2_NUM324_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM324 (.ZN (N1322), .A1 (XNOR_1_3_NAND2_NUM324_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM325_OUT, XNOR_1_2_NAND2_NUM325_OUT, XNOR_1_3_NAND2_NUM325_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM325 (.ZN (XNOR_1_1_NAND2_NUM325_OUT), .A1 (N730), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM325 (.ZN (XNOR_1_2_NAND2_NUM325_OUT), .A1 (GND), .A2 (N1238));
      NOR2_X1 XNOR_1_3_NAND2_NUM325 (.ZN (XNOR_1_3_NAND2_NUM325_OUT), .A1 (XNOR_1_1_NAND2_NUM325_OUT), .A2 (XNOR_1_2_NAND2_NUM325_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM325 (.ZN (N1327), .A1 (XNOR_1_3_NAND2_NUM325_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM326_OUT, XNOR_1_2_NAND2_NUM326_OUT, XNOR_1_3_NAND2_NUM326_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM326 (.ZN (XNOR_1_1_NAND2_NUM326_OUT), .A1 (N733), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM326 (.ZN (XNOR_1_2_NAND2_NUM326_OUT), .A1 (GND), .A2 (N1241));
      NOR2_X1 XNOR_1_3_NAND2_NUM326 (.ZN (XNOR_1_3_NAND2_NUM326_OUT), .A1 (XNOR_1_1_NAND2_NUM326_OUT), .A2 (XNOR_1_2_NAND2_NUM326_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM326 (.ZN (N1328), .A1 (XNOR_1_3_NAND2_NUM326_OUT), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM327 (.ZN (N1334), .A1 (N1162), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM328_OUT, XNOR_1_2_NAND2_NUM328_OUT, XNOR_1_3_NAND2_NUM328_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM328 (.ZN (XNOR_1_1_NAND2_NUM328_OUT), .A1 (N1267), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM328 (.ZN (XNOR_1_2_NAND2_NUM328_OUT), .A1 (GND), .A2 (N1160));
      NOR2_X1 XNOR_1_3_NAND2_NUM328 (.ZN (XNOR_1_3_NAND2_NUM328_OUT), .A1 (XNOR_1_1_NAND2_NUM328_OUT), .A2 (XNOR_1_2_NAND2_NUM328_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM328 (.ZN (N1344), .A1 (XNOR_1_3_NAND2_NUM328_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM329_OUT, XNOR_1_2_NAND2_NUM329_OUT, XNOR_1_3_NAND2_NUM329_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM329 (.ZN (XNOR_1_1_NAND2_NUM329_OUT), .A1 (N1249), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM329 (.ZN (XNOR_1_2_NAND2_NUM329_OUT), .A1 (GND), .A2 (N894));
      NOR2_X1 XNOR_1_3_NAND2_NUM329 (.ZN (XNOR_1_3_NAND2_NUM329_OUT), .A1 (XNOR_1_1_NAND2_NUM329_OUT), .A2 (XNOR_1_2_NAND2_NUM329_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM329 (.ZN (N1345), .A1 (XNOR_1_3_NAND2_NUM329_OUT), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM330 (.ZN (N1346), .A1 (N1249), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM331 (.ZN (N1348), .A1 (N1255), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM332 (.ZN (N1349), .A1 (N1252), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM333 (.ZN (N1350), .A1 (N1261), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM334 (.ZN (N1351), .A1 (N1258), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM335_OUT, XNOR_1_2_NAND2_NUM335_OUT, XNOR_1_3_NAND2_NUM335_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM335 (.ZN (XNOR_1_1_NAND2_NUM335_OUT), .A1 (N1309), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM335 (.ZN (XNOR_1_2_NAND2_NUM335_OUT), .A1 (GND), .A2 (N1206));
      NOR2_X1 XNOR_1_3_NAND2_NUM335 (.ZN (XNOR_1_3_NAND2_NUM335_OUT), .A1 (XNOR_1_1_NAND2_NUM335_OUT), .A2 (XNOR_1_2_NAND2_NUM335_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM335 (.ZN (N1352), .A1 (XNOR_1_3_NAND2_NUM335_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM336_OUT, XNOR_1_2_NAND2_NUM336_OUT, XNOR_1_3_NAND2_NUM336_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM336 (.ZN (XNOR_1_1_NAND2_NUM336_OUT), .A1 (N1310), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM336 (.ZN (XNOR_1_2_NAND2_NUM336_OUT), .A1 (GND), .A2 (N1208));
      NOR2_X1 XNOR_1_3_NAND2_NUM336 (.ZN (XNOR_1_3_NAND2_NUM336_OUT), .A1 (XNOR_1_1_NAND2_NUM336_OUT), .A2 (XNOR_1_2_NAND2_NUM336_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM336 (.ZN (N1355), .A1 (XNOR_1_3_NAND2_NUM336_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM337_OUT, XNOR_1_2_NAND2_NUM337_OUT, XNOR_1_3_NAND2_NUM337_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM337 (.ZN (XNOR_1_1_NAND2_NUM337_OUT), .A1 (N1311), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM337 (.ZN (XNOR_1_2_NAND2_NUM337_OUT), .A1 (GND), .A2 (N1210));
      NOR2_X1 XNOR_1_3_NAND2_NUM337 (.ZN (XNOR_1_3_NAND2_NUM337_OUT), .A1 (XNOR_1_1_NAND2_NUM337_OUT), .A2 (XNOR_1_2_NAND2_NUM337_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM337 (.ZN (N1358), .A1 (XNOR_1_3_NAND2_NUM337_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM338_OUT, XNOR_1_2_NAND2_NUM338_OUT, XNOR_1_3_NAND2_NUM338_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM338 (.ZN (XNOR_1_1_NAND2_NUM338_OUT), .A1 (N1312), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM338 (.ZN (XNOR_1_2_NAND2_NUM338_OUT), .A1 (GND), .A2 (N1212));
      NOR2_X1 XNOR_1_3_NAND2_NUM338 (.ZN (XNOR_1_3_NAND2_NUM338_OUT), .A1 (XNOR_1_1_NAND2_NUM338_OUT), .A2 (XNOR_1_2_NAND2_NUM338_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM338 (.ZN (N1361), .A1 (XNOR_1_3_NAND2_NUM338_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM339_OUT, XNOR_1_2_NAND2_NUM339_OUT, XNOR_1_3_NAND2_NUM339_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM339 (.ZN (XNOR_1_1_NAND2_NUM339_OUT), .A1 (N1313), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM339 (.ZN (XNOR_1_2_NAND2_NUM339_OUT), .A1 (GND), .A2 (N1214));
      NOR2_X1 XNOR_1_3_NAND2_NUM339 (.ZN (XNOR_1_3_NAND2_NUM339_OUT), .A1 (XNOR_1_1_NAND2_NUM339_OUT), .A2 (XNOR_1_2_NAND2_NUM339_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM339 (.ZN (N1364), .A1 (XNOR_1_3_NAND2_NUM339_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM340_OUT, XNOR_1_2_NAND2_NUM340_OUT, XNOR_1_3_NAND2_NUM340_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM340 (.ZN (XNOR_1_1_NAND2_NUM340_OUT), .A1 (N1314), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM340 (.ZN (XNOR_1_2_NAND2_NUM340_OUT), .A1 (GND), .A2 (N1216));
      NOR2_X1 XNOR_1_3_NAND2_NUM340 (.ZN (XNOR_1_3_NAND2_NUM340_OUT), .A1 (XNOR_1_1_NAND2_NUM340_OUT), .A2 (XNOR_1_2_NAND2_NUM340_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM340 (.ZN (N1367), .A1 (XNOR_1_3_NAND2_NUM340_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM341_OUT, XNOR_1_2_NAND2_NUM341_OUT, XNOR_1_3_NAND2_NUM341_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM341 (.ZN (XNOR_1_1_NAND2_NUM341_OUT), .A1 (N1315), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM341 (.ZN (XNOR_1_2_NAND2_NUM341_OUT), .A1 (GND), .A2 (N1221));
      NOR2_X1 XNOR_1_3_NAND2_NUM341 (.ZN (XNOR_1_3_NAND2_NUM341_OUT), .A1 (XNOR_1_1_NAND2_NUM341_OUT), .A2 (XNOR_1_2_NAND2_NUM341_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM341 (.ZN (N1370), .A1 (XNOR_1_3_NAND2_NUM341_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM342_OUT, XNOR_1_2_NAND2_NUM342_OUT, XNOR_1_3_NAND2_NUM342_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM342 (.ZN (XNOR_1_1_NAND2_NUM342_OUT), .A1 (N1316), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM342 (.ZN (XNOR_1_2_NAND2_NUM342_OUT), .A1 (GND), .A2 (N1224));
      NOR2_X1 XNOR_1_3_NAND2_NUM342 (.ZN (XNOR_1_3_NAND2_NUM342_OUT), .A1 (XNOR_1_1_NAND2_NUM342_OUT), .A2 (XNOR_1_2_NAND2_NUM342_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM342 (.ZN (N1373), .A1 (XNOR_1_3_NAND2_NUM342_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM343_OUT, XNOR_1_2_NAND2_NUM343_OUT, XNOR_1_3_NAND2_NUM343_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM343 (.ZN (XNOR_1_1_NAND2_NUM343_OUT), .A1 (N1317), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM343 (.ZN (XNOR_1_2_NAND2_NUM343_OUT), .A1 (GND), .A2 (N1226));
      NOR2_X1 XNOR_1_3_NAND2_NUM343 (.ZN (XNOR_1_3_NAND2_NUM343_OUT), .A1 (XNOR_1_1_NAND2_NUM343_OUT), .A2 (XNOR_1_2_NAND2_NUM343_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM343 (.ZN (N1376), .A1 (XNOR_1_3_NAND2_NUM343_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM344_OUT, XNOR_1_2_NAND2_NUM344_OUT, XNOR_1_3_NAND2_NUM344_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM344 (.ZN (XNOR_1_1_NAND2_NUM344_OUT), .A1 (N1318), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM344 (.ZN (XNOR_1_2_NAND2_NUM344_OUT), .A1 (GND), .A2 (N1229));
      NOR2_X1 XNOR_1_3_NAND2_NUM344 (.ZN (XNOR_1_3_NAND2_NUM344_OUT), .A1 (XNOR_1_1_NAND2_NUM344_OUT), .A2 (XNOR_1_2_NAND2_NUM344_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM344 (.ZN (N1379), .A1 (XNOR_1_3_NAND2_NUM344_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM345_OUT, XNOR_1_2_NAND2_NUM345_OUT, XNOR_1_3_NAND2_NUM345_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM345 (.ZN (XNOR_1_1_NAND2_NUM345_OUT), .A1 (N1322), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM345 (.ZN (XNOR_1_2_NAND2_NUM345_OUT), .A1 (GND), .A2 (N1231));
      NOR2_X1 XNOR_1_3_NAND2_NUM345 (.ZN (XNOR_1_3_NAND2_NUM345_OUT), .A1 (XNOR_1_1_NAND2_NUM345_OUT), .A2 (XNOR_1_2_NAND2_NUM345_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM345 (.ZN (N1383), .A1 (XNOR_1_3_NAND2_NUM345_OUT), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM346 (.ZN (N1386), .A1 (N1232), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM347_OUT, XNOR_1_2_NAND2_NUM347_OUT, XNOR_1_3_NAND2_NUM347_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM347 (.ZN (XNOR_1_1_NAND2_NUM347_OUT), .A1 (N1232), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM347 (.ZN (XNOR_1_2_NAND2_NUM347_OUT), .A1 (GND), .A2 (N990));
      NOR2_X1 XNOR_1_3_NAND2_NUM347 (.ZN (XNOR_1_3_NAND2_NUM347_OUT), .A1 (XNOR_1_1_NAND2_NUM347_OUT), .A2 (XNOR_1_2_NAND2_NUM347_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM347 (.ZN (N1387), .A1 (XNOR_1_3_NAND2_NUM347_OUT), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM348 (.ZN (N1388), .A1 (N1235), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM349_OUT, XNOR_1_2_NAND2_NUM349_OUT, XNOR_1_3_NAND2_NUM349_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM349 (.ZN (XNOR_1_1_NAND2_NUM349_OUT), .A1 (N1235), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM349 (.ZN (XNOR_1_2_NAND2_NUM349_OUT), .A1 (GND), .A2 (N993));
      NOR2_X1 XNOR_1_3_NAND2_NUM349 (.ZN (XNOR_1_3_NAND2_NUM349_OUT), .A1 (XNOR_1_1_NAND2_NUM349_OUT), .A2 (XNOR_1_2_NAND2_NUM349_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM349 (.ZN (N1389), .A1 (XNOR_1_3_NAND2_NUM349_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM350_OUT, XNOR_1_2_NAND2_NUM350_OUT, XNOR_1_3_NAND2_NUM350_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM350 (.ZN (XNOR_1_1_NAND2_NUM350_OUT), .A1 (N1327), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM350 (.ZN (XNOR_1_2_NAND2_NUM350_OUT), .A1 (GND), .A2 (N1239));
      NOR2_X1 XNOR_1_3_NAND2_NUM350 (.ZN (XNOR_1_3_NAND2_NUM350_OUT), .A1 (XNOR_1_1_NAND2_NUM350_OUT), .A2 (XNOR_1_2_NAND2_NUM350_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM350 (.ZN (N1390), .A1 (XNOR_1_3_NAND2_NUM350_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM351_OUT, XNOR_1_2_NAND2_NUM351_OUT, XNOR_1_3_NAND2_NUM351_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM351 (.ZN (XNOR_1_1_NAND2_NUM351_OUT), .A1 (N1328), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM351 (.ZN (XNOR_1_2_NAND2_NUM351_OUT), .A1 (GND), .A2 (N1242));
      NOR2_X1 XNOR_1_3_NAND2_NUM351 (.ZN (XNOR_1_3_NAND2_NUM351_OUT), .A1 (XNOR_1_1_NAND2_NUM351_OUT), .A2 (XNOR_1_2_NAND2_NUM351_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM351 (.ZN (N1393), .A1 (XNOR_1_3_NAND2_NUM351_OUT), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM352 (.ZN (N1396), .A1 (N1243), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM353_OUT, XNOR_1_2_NAND2_NUM353_OUT, XNOR_1_3_NAND2_NUM353_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM353 (.ZN (XNOR_1_1_NAND2_NUM353_OUT), .A1 (N1243), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM353 (.ZN (XNOR_1_2_NAND2_NUM353_OUT), .A1 (GND), .A2 (N1004));
      NOR2_X1 XNOR_1_3_NAND2_NUM353 (.ZN (XNOR_1_3_NAND2_NUM353_OUT), .A1 (XNOR_1_1_NAND2_NUM353_OUT), .A2 (XNOR_1_2_NAND2_NUM353_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM353 (.ZN (N1397), .A1 (XNOR_1_3_NAND2_NUM353_OUT), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM354 (.ZN (N1398), .A1 (N1246), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM355_OUT, XNOR_1_2_NAND2_NUM355_OUT, XNOR_1_3_NAND2_NUM355_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM355 (.ZN (XNOR_1_1_NAND2_NUM355_OUT), .A1 (N1246), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM355 (.ZN (XNOR_1_2_NAND2_NUM355_OUT), .A1 (GND), .A2 (N1007));
      NOR2_X1 XNOR_1_3_NAND2_NUM355 (.ZN (XNOR_1_3_NAND2_NUM355_OUT), .A1 (XNOR_1_1_NAND2_NUM355_OUT), .A2 (XNOR_1_2_NAND2_NUM355_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM355 (.ZN (N1399), .A1 (XNOR_1_3_NAND2_NUM355_OUT), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM356 (.ZN (N1409), .A1 (N1319), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM357_OUT, XNOR_1_2_NAND2_NUM357_OUT, XNOR_1_3_NAND2_NUM357_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM357 (.ZN (XNOR_1_1_NAND2_NUM357_OUT), .A1 (N649), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM357 (.ZN (XNOR_1_2_NAND2_NUM357_OUT), .A1 (GND), .A2 (N1346));
      NOR2_X1 XNOR_1_3_NAND2_NUM357 (.ZN (XNOR_1_3_NAND2_NUM357_OUT), .A1 (XNOR_1_1_NAND2_NUM357_OUT), .A2 (XNOR_1_2_NAND2_NUM357_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM357 (.ZN (N1412), .A1 (XNOR_1_3_NAND2_NUM357_OUT), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM358 (.ZN (N1413), .A1 (N1334), .A2 (GND));
      wire XNOR_1_1_BUFF1_NUM359_OUT;
      NOR2_X1 XNOR_1_1_BUFF1_NUM359 (.ZN (XNOR_1_1_BUFF1_NUM359_OUT), .A1 (N1264), .A2 (GND));
      NOR2_X1 XNOR_1_2_BUFF1_NUM359 (.ZN (N1416), .A1 (XNOR_1_1_BUFF1_NUM359_OUT), .A2 (GND));
      wire XNOR_1_1_BUFF1_NUM360_OUT;
      NOR2_X1 XNOR_1_1_BUFF1_NUM360 (.ZN (XNOR_1_1_BUFF1_NUM360_OUT), .A1 (N1264), .A2 (GND));
      NOR2_X1 XNOR_1_2_BUFF1_NUM360 (.ZN (N1419), .A1 (XNOR_1_1_BUFF1_NUM360_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM361_OUT, XNOR_1_2_NAND2_NUM361_OUT, XNOR_1_3_NAND2_NUM361_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM361 (.ZN (XNOR_1_1_NAND2_NUM361_OUT), .A1 (N634), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM361 (.ZN (XNOR_1_2_NAND2_NUM361_OUT), .A1 (GND), .A2 (N1386));
      NOR2_X1 XNOR_1_3_NAND2_NUM361 (.ZN (XNOR_1_3_NAND2_NUM361_OUT), .A1 (XNOR_1_1_NAND2_NUM361_OUT), .A2 (XNOR_1_2_NAND2_NUM361_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM361 (.ZN (N1433), .A1 (XNOR_1_3_NAND2_NUM361_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM362_OUT, XNOR_1_2_NAND2_NUM362_OUT, XNOR_1_3_NAND2_NUM362_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM362 (.ZN (XNOR_1_1_NAND2_NUM362_OUT), .A1 (N637), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM362 (.ZN (XNOR_1_2_NAND2_NUM362_OUT), .A1 (GND), .A2 (N1388));
      NOR2_X1 XNOR_1_3_NAND2_NUM362 (.ZN (XNOR_1_3_NAND2_NUM362_OUT), .A1 (XNOR_1_1_NAND2_NUM362_OUT), .A2 (XNOR_1_2_NAND2_NUM362_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM362 (.ZN (N1434), .A1 (XNOR_1_3_NAND2_NUM362_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM363_OUT, XNOR_1_2_NAND2_NUM363_OUT, XNOR_1_3_NAND2_NUM363_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM363 (.ZN (XNOR_1_1_NAND2_NUM363_OUT), .A1 (N640), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM363 (.ZN (XNOR_1_2_NAND2_NUM363_OUT), .A1 (GND), .A2 (N1396));
      NOR2_X1 XNOR_1_3_NAND2_NUM363 (.ZN (XNOR_1_3_NAND2_NUM363_OUT), .A1 (XNOR_1_1_NAND2_NUM363_OUT), .A2 (XNOR_1_2_NAND2_NUM363_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM363 (.ZN (N1438), .A1 (XNOR_1_3_NAND2_NUM363_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM364_OUT, XNOR_1_2_NAND2_NUM364_OUT, XNOR_1_3_NAND2_NUM364_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM364 (.ZN (XNOR_1_1_NAND2_NUM364_OUT), .A1 (N646), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM364 (.ZN (XNOR_1_2_NAND2_NUM364_OUT), .A1 (GND), .A2 (N1398));
      NOR2_X1 XNOR_1_3_NAND2_NUM364 (.ZN (XNOR_1_3_NAND2_NUM364_OUT), .A1 (XNOR_1_1_NAND2_NUM364_OUT), .A2 (XNOR_1_2_NAND2_NUM364_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM364 (.ZN (N1439), .A1 (XNOR_1_3_NAND2_NUM364_OUT), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM365 (.ZN (N1440), .A1 (N1344), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM366_OUT, XNOR_1_2_NAND2_NUM366_OUT, XNOR_1_3_NAND2_NUM366_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM366 (.ZN (XNOR_1_1_NAND2_NUM366_OUT), .A1 (N1355), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM366 (.ZN (XNOR_1_2_NAND2_NUM366_OUT), .A1 (GND), .A2 (N1148));
      NOR2_X1 XNOR_1_3_NAND2_NUM366 (.ZN (XNOR_1_3_NAND2_NUM366_OUT), .A1 (XNOR_1_1_NAND2_NUM366_OUT), .A2 (XNOR_1_2_NAND2_NUM366_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM366 (.ZN (N1443), .A1 (XNOR_1_3_NAND2_NUM366_OUT), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM367 (.ZN (N1444), .A1 (N1355), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM368_OUT, XNOR_1_2_NAND2_NUM368_OUT, XNOR_1_3_NAND2_NUM368_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM368 (.ZN (XNOR_1_1_NAND2_NUM368_OUT), .A1 (N1352), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM368 (.ZN (XNOR_1_2_NAND2_NUM368_OUT), .A1 (GND), .A2 (N1149));
      NOR2_X1 XNOR_1_3_NAND2_NUM368 (.ZN (XNOR_1_3_NAND2_NUM368_OUT), .A1 (XNOR_1_1_NAND2_NUM368_OUT), .A2 (XNOR_1_2_NAND2_NUM368_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM368 (.ZN (N1445), .A1 (XNOR_1_3_NAND2_NUM368_OUT), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM369 (.ZN (N1446), .A1 (N1352), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM370_OUT, XNOR_1_2_NAND2_NUM370_OUT, XNOR_1_3_NAND2_NUM370_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM370 (.ZN (XNOR_1_1_NAND2_NUM370_OUT), .A1 (N1358), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM370 (.ZN (XNOR_1_2_NAND2_NUM370_OUT), .A1 (GND), .A2 (N1151));
      NOR2_X1 XNOR_1_3_NAND2_NUM370 (.ZN (XNOR_1_3_NAND2_NUM370_OUT), .A1 (XNOR_1_1_NAND2_NUM370_OUT), .A2 (XNOR_1_2_NAND2_NUM370_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM370 (.ZN (N1447), .A1 (XNOR_1_3_NAND2_NUM370_OUT), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM371 (.ZN (N1448), .A1 (N1358), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM372_OUT, XNOR_1_2_NAND2_NUM372_OUT, XNOR_1_3_NAND2_NUM372_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM372 (.ZN (XNOR_1_1_NAND2_NUM372_OUT), .A1 (N1361), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM372 (.ZN (XNOR_1_2_NAND2_NUM372_OUT), .A1 (GND), .A2 (N1152));
      NOR2_X1 XNOR_1_3_NAND2_NUM372 (.ZN (XNOR_1_3_NAND2_NUM372_OUT), .A1 (XNOR_1_1_NAND2_NUM372_OUT), .A2 (XNOR_1_2_NAND2_NUM372_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM372 (.ZN (N1451), .A1 (XNOR_1_3_NAND2_NUM372_OUT), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM373 (.ZN (N1452), .A1 (N1361), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM374_OUT, XNOR_1_2_NAND2_NUM374_OUT, XNOR_1_3_NAND2_NUM374_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM374 (.ZN (XNOR_1_1_NAND2_NUM374_OUT), .A1 (N1367), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM374 (.ZN (XNOR_1_2_NAND2_NUM374_OUT), .A1 (GND), .A2 (N1153));
      NOR2_X1 XNOR_1_3_NAND2_NUM374 (.ZN (XNOR_1_3_NAND2_NUM374_OUT), .A1 (XNOR_1_1_NAND2_NUM374_OUT), .A2 (XNOR_1_2_NAND2_NUM374_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM374 (.ZN (N1453), .A1 (XNOR_1_3_NAND2_NUM374_OUT), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM375 (.ZN (N1454), .A1 (N1367), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM376_OUT, XNOR_1_2_NAND2_NUM376_OUT, XNOR_1_3_NAND2_NUM376_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM376 (.ZN (XNOR_1_1_NAND2_NUM376_OUT), .A1 (N1364), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM376 (.ZN (XNOR_1_2_NAND2_NUM376_OUT), .A1 (GND), .A2 (N1154));
      NOR2_X1 XNOR_1_3_NAND2_NUM376 (.ZN (XNOR_1_3_NAND2_NUM376_OUT), .A1 (XNOR_1_1_NAND2_NUM376_OUT), .A2 (XNOR_1_2_NAND2_NUM376_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM376 (.ZN (N1455), .A1 (XNOR_1_3_NAND2_NUM376_OUT), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM377 (.ZN (N1456), .A1 (N1364), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM378_OUT, XNOR_1_2_NAND2_NUM378_OUT, XNOR_1_3_NAND2_NUM378_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM378 (.ZN (XNOR_1_1_NAND2_NUM378_OUT), .A1 (N1373), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM378 (.ZN (XNOR_1_2_NAND2_NUM378_OUT), .A1 (GND), .A2 (N1156));
      NOR2_X1 XNOR_1_3_NAND2_NUM378 (.ZN (XNOR_1_3_NAND2_NUM378_OUT), .A1 (XNOR_1_1_NAND2_NUM378_OUT), .A2 (XNOR_1_2_NAND2_NUM378_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM378 (.ZN (N1457), .A1 (XNOR_1_3_NAND2_NUM378_OUT), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM379 (.ZN (N1458), .A1 (N1373), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM380_OUT, XNOR_1_2_NAND2_NUM380_OUT, XNOR_1_3_NAND2_NUM380_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM380 (.ZN (XNOR_1_1_NAND2_NUM380_OUT), .A1 (N1379), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM380 (.ZN (XNOR_1_2_NAND2_NUM380_OUT), .A1 (GND), .A2 (N1157));
      NOR2_X1 XNOR_1_3_NAND2_NUM380 (.ZN (XNOR_1_3_NAND2_NUM380_OUT), .A1 (XNOR_1_1_NAND2_NUM380_OUT), .A2 (XNOR_1_2_NAND2_NUM380_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM380 (.ZN (N1459), .A1 (XNOR_1_3_NAND2_NUM380_OUT), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM381 (.ZN (N1460), .A1 (N1379), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM382 (.ZN (N1461), .A1 (N1383), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM383_OUT, XNOR_1_2_NAND2_NUM383_OUT, XNOR_1_3_NAND2_NUM383_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM383 (.ZN (XNOR_1_1_NAND2_NUM383_OUT), .A1 (N1393), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM383 (.ZN (XNOR_1_2_NAND2_NUM383_OUT), .A1 (GND), .A2 (N1161));
      NOR2_X1 XNOR_1_3_NAND2_NUM383 (.ZN (XNOR_1_3_NAND2_NUM383_OUT), .A1 (XNOR_1_1_NAND2_NUM383_OUT), .A2 (XNOR_1_2_NAND2_NUM383_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM383 (.ZN (N1462), .A1 (XNOR_1_3_NAND2_NUM383_OUT), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM384 (.ZN (N1463), .A1 (N1393), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM385_OUT, XNOR_1_2_NAND2_NUM385_OUT, XNOR_1_3_NAND2_NUM385_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM385 (.ZN (XNOR_1_1_NAND2_NUM385_OUT), .A1 (N1345), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM385 (.ZN (XNOR_1_2_NAND2_NUM385_OUT), .A1 (GND), .A2 (N1412));
      NOR2_X1 XNOR_1_3_NAND2_NUM385 (.ZN (XNOR_1_3_NAND2_NUM385_OUT), .A1 (XNOR_1_1_NAND2_NUM385_OUT), .A2 (XNOR_1_2_NAND2_NUM385_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM385 (.ZN (N1464), .A1 (XNOR_1_3_NAND2_NUM385_OUT), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM386 (.ZN (N1468), .A1 (N1370), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM387_OUT, XNOR_1_2_NAND2_NUM387_OUT, XNOR_1_3_NAND2_NUM387_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM387 (.ZN (XNOR_1_1_NAND2_NUM387_OUT), .A1 (N1370), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM387 (.ZN (XNOR_1_2_NAND2_NUM387_OUT), .A1 (GND), .A2 (N1222));
      NOR2_X1 XNOR_1_3_NAND2_NUM387 (.ZN (XNOR_1_3_NAND2_NUM387_OUT), .A1 (XNOR_1_1_NAND2_NUM387_OUT), .A2 (XNOR_1_2_NAND2_NUM387_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM387 (.ZN (N1469), .A1 (XNOR_1_3_NAND2_NUM387_OUT), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM388 (.ZN (N1470), .A1 (N1376), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM389_OUT, XNOR_1_2_NAND2_NUM389_OUT, XNOR_1_3_NAND2_NUM389_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM389 (.ZN (XNOR_1_1_NAND2_NUM389_OUT), .A1 (N1376), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM389 (.ZN (XNOR_1_2_NAND2_NUM389_OUT), .A1 (GND), .A2 (N1227));
      NOR2_X1 XNOR_1_3_NAND2_NUM389 (.ZN (XNOR_1_3_NAND2_NUM389_OUT), .A1 (XNOR_1_1_NAND2_NUM389_OUT), .A2 (XNOR_1_2_NAND2_NUM389_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM389 (.ZN (N1471), .A1 (XNOR_1_3_NAND2_NUM389_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM390_OUT, XNOR_1_2_NAND2_NUM390_OUT, XNOR_1_3_NAND2_NUM390_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM390 (.ZN (XNOR_1_1_NAND2_NUM390_OUT), .A1 (N1387), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM390 (.ZN (XNOR_1_2_NAND2_NUM390_OUT), .A1 (GND), .A2 (N1433));
      NOR2_X1 XNOR_1_3_NAND2_NUM390 (.ZN (XNOR_1_3_NAND2_NUM390_OUT), .A1 (XNOR_1_1_NAND2_NUM390_OUT), .A2 (XNOR_1_2_NAND2_NUM390_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM390 (.ZN (N1472), .A1 (XNOR_1_3_NAND2_NUM390_OUT), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM391 (.ZN (N1475), .A1 (N1390), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM392_OUT, XNOR_1_2_NAND2_NUM392_OUT, XNOR_1_3_NAND2_NUM392_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM392 (.ZN (XNOR_1_1_NAND2_NUM392_OUT), .A1 (N1390), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM392 (.ZN (XNOR_1_2_NAND2_NUM392_OUT), .A1 (GND), .A2 (N1240));
      NOR2_X1 XNOR_1_3_NAND2_NUM392 (.ZN (XNOR_1_3_NAND2_NUM392_OUT), .A1 (XNOR_1_1_NAND2_NUM392_OUT), .A2 (XNOR_1_2_NAND2_NUM392_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM392 (.ZN (N1476), .A1 (XNOR_1_3_NAND2_NUM392_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM393_OUT, XNOR_1_2_NAND2_NUM393_OUT, XNOR_1_3_NAND2_NUM393_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM393 (.ZN (XNOR_1_1_NAND2_NUM393_OUT), .A1 (N1389), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM393 (.ZN (XNOR_1_2_NAND2_NUM393_OUT), .A1 (GND), .A2 (N1434));
      NOR2_X1 XNOR_1_3_NAND2_NUM393 (.ZN (XNOR_1_3_NAND2_NUM393_OUT), .A1 (XNOR_1_1_NAND2_NUM393_OUT), .A2 (XNOR_1_2_NAND2_NUM393_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM393 (.ZN (N1478), .A1 (XNOR_1_3_NAND2_NUM393_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM394_OUT, XNOR_1_2_NAND2_NUM394_OUT, XNOR_1_3_NAND2_NUM394_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM394 (.ZN (XNOR_1_1_NAND2_NUM394_OUT), .A1 (N1399), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM394 (.ZN (XNOR_1_2_NAND2_NUM394_OUT), .A1 (GND), .A2 (N1439));
      NOR2_X1 XNOR_1_3_NAND2_NUM394 (.ZN (XNOR_1_3_NAND2_NUM394_OUT), .A1 (XNOR_1_1_NAND2_NUM394_OUT), .A2 (XNOR_1_2_NAND2_NUM394_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM394 (.ZN (N1481), .A1 (XNOR_1_3_NAND2_NUM394_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM395_OUT, XNOR_1_2_NAND2_NUM395_OUT, XNOR_1_3_NAND2_NUM395_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM395 (.ZN (XNOR_1_1_NAND2_NUM395_OUT), .A1 (N1397), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM395 (.ZN (XNOR_1_2_NAND2_NUM395_OUT), .A1 (GND), .A2 (N1438));
      NOR2_X1 XNOR_1_3_NAND2_NUM395 (.ZN (XNOR_1_3_NAND2_NUM395_OUT), .A1 (XNOR_1_1_NAND2_NUM395_OUT), .A2 (XNOR_1_2_NAND2_NUM395_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM395 (.ZN (N1484), .A1 (XNOR_1_3_NAND2_NUM395_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM396_OUT, XNOR_1_2_NAND2_NUM396_OUT, XNOR_1_3_NAND2_NUM396_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM396 (.ZN (XNOR_1_1_NAND2_NUM396_OUT), .A1 (N939), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM396 (.ZN (XNOR_1_2_NAND2_NUM396_OUT), .A1 (GND), .A2 (N1444));
      NOR2_X1 XNOR_1_3_NAND2_NUM396 (.ZN (XNOR_1_3_NAND2_NUM396_OUT), .A1 (XNOR_1_1_NAND2_NUM396_OUT), .A2 (XNOR_1_2_NAND2_NUM396_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM396 (.ZN (N1487), .A1 (XNOR_1_3_NAND2_NUM396_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM397_OUT, XNOR_1_2_NAND2_NUM397_OUT, XNOR_1_3_NAND2_NUM397_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM397 (.ZN (XNOR_1_1_NAND2_NUM397_OUT), .A1 (N935), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM397 (.ZN (XNOR_1_2_NAND2_NUM397_OUT), .A1 (GND), .A2 (N1446));
      NOR2_X1 XNOR_1_3_NAND2_NUM397 (.ZN (XNOR_1_3_NAND2_NUM397_OUT), .A1 (XNOR_1_1_NAND2_NUM397_OUT), .A2 (XNOR_1_2_NAND2_NUM397_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM397 (.ZN (N1488), .A1 (XNOR_1_3_NAND2_NUM397_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM398_OUT, XNOR_1_2_NAND2_NUM398_OUT, XNOR_1_3_NAND2_NUM398_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM398 (.ZN (XNOR_1_1_NAND2_NUM398_OUT), .A1 (N943), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM398 (.ZN (XNOR_1_2_NAND2_NUM398_OUT), .A1 (GND), .A2 (N1448));
      NOR2_X1 XNOR_1_3_NAND2_NUM398 (.ZN (XNOR_1_3_NAND2_NUM398_OUT), .A1 (XNOR_1_1_NAND2_NUM398_OUT), .A2 (XNOR_1_2_NAND2_NUM398_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM398 (.ZN (N1489), .A1 (XNOR_1_3_NAND2_NUM398_OUT), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM399 (.ZN (N1490), .A1 (N1419), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM400 (.ZN (N1491), .A1 (N1416), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM401_OUT, XNOR_1_2_NAND2_NUM401_OUT, XNOR_1_3_NAND2_NUM401_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM401 (.ZN (XNOR_1_1_NAND2_NUM401_OUT), .A1 (N947), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM401 (.ZN (XNOR_1_2_NAND2_NUM401_OUT), .A1 (GND), .A2 (N1452));
      NOR2_X1 XNOR_1_3_NAND2_NUM401 (.ZN (XNOR_1_3_NAND2_NUM401_OUT), .A1 (XNOR_1_1_NAND2_NUM401_OUT), .A2 (XNOR_1_2_NAND2_NUM401_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM401 (.ZN (N1492), .A1 (XNOR_1_3_NAND2_NUM401_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM402_OUT, XNOR_1_2_NAND2_NUM402_OUT, XNOR_1_3_NAND2_NUM402_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM402 (.ZN (XNOR_1_1_NAND2_NUM402_OUT), .A1 (N955), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM402 (.ZN (XNOR_1_2_NAND2_NUM402_OUT), .A1 (GND), .A2 (N1454));
      NOR2_X1 XNOR_1_3_NAND2_NUM402 (.ZN (XNOR_1_3_NAND2_NUM402_OUT), .A1 (XNOR_1_1_NAND2_NUM402_OUT), .A2 (XNOR_1_2_NAND2_NUM402_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM402 (.ZN (N1493), .A1 (XNOR_1_3_NAND2_NUM402_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM403_OUT, XNOR_1_2_NAND2_NUM403_OUT, XNOR_1_3_NAND2_NUM403_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM403 (.ZN (XNOR_1_1_NAND2_NUM403_OUT), .A1 (N951), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM403 (.ZN (XNOR_1_2_NAND2_NUM403_OUT), .A1 (GND), .A2 (N1456));
      NOR2_X1 XNOR_1_3_NAND2_NUM403 (.ZN (XNOR_1_3_NAND2_NUM403_OUT), .A1 (XNOR_1_1_NAND2_NUM403_OUT), .A2 (XNOR_1_2_NAND2_NUM403_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM403 (.ZN (N1494), .A1 (XNOR_1_3_NAND2_NUM403_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM404_OUT, XNOR_1_2_NAND2_NUM404_OUT, XNOR_1_3_NAND2_NUM404_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM404 (.ZN (XNOR_1_1_NAND2_NUM404_OUT), .A1 (N969), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM404 (.ZN (XNOR_1_2_NAND2_NUM404_OUT), .A1 (GND), .A2 (N1458));
      NOR2_X1 XNOR_1_3_NAND2_NUM404 (.ZN (XNOR_1_3_NAND2_NUM404_OUT), .A1 (XNOR_1_1_NAND2_NUM404_OUT), .A2 (XNOR_1_2_NAND2_NUM404_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM404 (.ZN (N1495), .A1 (XNOR_1_3_NAND2_NUM404_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM405_OUT, XNOR_1_2_NAND2_NUM405_OUT, XNOR_1_3_NAND2_NUM405_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM405 (.ZN (XNOR_1_1_NAND2_NUM405_OUT), .A1 (N977), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM405 (.ZN (XNOR_1_2_NAND2_NUM405_OUT), .A1 (GND), .A2 (N1460));
      NOR2_X1 XNOR_1_3_NAND2_NUM405 (.ZN (XNOR_1_3_NAND2_NUM405_OUT), .A1 (XNOR_1_1_NAND2_NUM405_OUT), .A2 (XNOR_1_2_NAND2_NUM405_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM405 (.ZN (N1496), .A1 (XNOR_1_3_NAND2_NUM405_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM406_OUT, XNOR_1_2_NAND2_NUM406_OUT, XNOR_1_3_NAND2_NUM406_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM406 (.ZN (XNOR_1_1_NAND2_NUM406_OUT), .A1 (N998), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM406 (.ZN (XNOR_1_2_NAND2_NUM406_OUT), .A1 (GND), .A2 (N1463));
      NOR2_X1 XNOR_1_3_NAND2_NUM406 (.ZN (XNOR_1_3_NAND2_NUM406_OUT), .A1 (XNOR_1_1_NAND2_NUM406_OUT), .A2 (XNOR_1_2_NAND2_NUM406_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM406 (.ZN (N1498), .A1 (XNOR_1_3_NAND2_NUM406_OUT), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM407 (.ZN (N1499), .A1 (N1440), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM408_OUT, XNOR_1_2_NAND2_NUM408_OUT, XNOR_1_3_NAND2_NUM408_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM408 (.ZN (XNOR_1_1_NAND2_NUM408_OUT), .A1 (N965), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM408 (.ZN (XNOR_1_2_NAND2_NUM408_OUT), .A1 (GND), .A2 (N1468));
      NOR2_X1 XNOR_1_3_NAND2_NUM408 (.ZN (XNOR_1_3_NAND2_NUM408_OUT), .A1 (XNOR_1_1_NAND2_NUM408_OUT), .A2 (XNOR_1_2_NAND2_NUM408_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM408 (.ZN (N1500), .A1 (XNOR_1_3_NAND2_NUM408_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM409_OUT, XNOR_1_2_NAND2_NUM409_OUT, XNOR_1_3_NAND2_NUM409_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM409 (.ZN (XNOR_1_1_NAND2_NUM409_OUT), .A1 (N973), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM409 (.ZN (XNOR_1_2_NAND2_NUM409_OUT), .A1 (GND), .A2 (N1470));
      NOR2_X1 XNOR_1_3_NAND2_NUM409 (.ZN (XNOR_1_3_NAND2_NUM409_OUT), .A1 (XNOR_1_1_NAND2_NUM409_OUT), .A2 (XNOR_1_2_NAND2_NUM409_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM409 (.ZN (N1501), .A1 (XNOR_1_3_NAND2_NUM409_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM410_OUT, XNOR_1_2_NAND2_NUM410_OUT, XNOR_1_3_NAND2_NUM410_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM410 (.ZN (XNOR_1_1_NAND2_NUM410_OUT), .A1 (N994), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM410 (.ZN (XNOR_1_2_NAND2_NUM410_OUT), .A1 (GND), .A2 (N1475));
      NOR2_X1 XNOR_1_3_NAND2_NUM410 (.ZN (XNOR_1_3_NAND2_NUM410_OUT), .A1 (XNOR_1_1_NAND2_NUM410_OUT), .A2 (XNOR_1_2_NAND2_NUM410_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM410 (.ZN (N1504), .A1 (XNOR_1_3_NAND2_NUM410_OUT), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM411 (.ZN (N1510), .A1 (N1464), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM412_OUT, XNOR_1_2_NAND2_NUM412_OUT, XNOR_1_3_NAND2_NUM412_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM412 (.ZN (XNOR_1_1_NAND2_NUM412_OUT), .A1 (N1443), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM412 (.ZN (XNOR_1_2_NAND2_NUM412_OUT), .A1 (GND), .A2 (N1487));
      NOR2_X1 XNOR_1_3_NAND2_NUM412 (.ZN (XNOR_1_3_NAND2_NUM412_OUT), .A1 (XNOR_1_1_NAND2_NUM412_OUT), .A2 (XNOR_1_2_NAND2_NUM412_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM412 (.ZN (N1513), .A1 (XNOR_1_3_NAND2_NUM412_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM413_OUT, XNOR_1_2_NAND2_NUM413_OUT, XNOR_1_3_NAND2_NUM413_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM413 (.ZN (XNOR_1_1_NAND2_NUM413_OUT), .A1 (N1445), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM413 (.ZN (XNOR_1_2_NAND2_NUM413_OUT), .A1 (GND), .A2 (N1488));
      NOR2_X1 XNOR_1_3_NAND2_NUM413 (.ZN (XNOR_1_3_NAND2_NUM413_OUT), .A1 (XNOR_1_1_NAND2_NUM413_OUT), .A2 (XNOR_1_2_NAND2_NUM413_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM413 (.ZN (N1514), .A1 (XNOR_1_3_NAND2_NUM413_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM414_OUT, XNOR_1_2_NAND2_NUM414_OUT, XNOR_1_3_NAND2_NUM414_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM414 (.ZN (XNOR_1_1_NAND2_NUM414_OUT), .A1 (N1447), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM414 (.ZN (XNOR_1_2_NAND2_NUM414_OUT), .A1 (GND), .A2 (N1489));
      NOR2_X1 XNOR_1_3_NAND2_NUM414 (.ZN (XNOR_1_3_NAND2_NUM414_OUT), .A1 (XNOR_1_1_NAND2_NUM414_OUT), .A2 (XNOR_1_2_NAND2_NUM414_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM414 (.ZN (N1517), .A1 (XNOR_1_3_NAND2_NUM414_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM415_OUT, XNOR_1_2_NAND2_NUM415_OUT, XNOR_1_3_NAND2_NUM415_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM415 (.ZN (XNOR_1_1_NAND2_NUM415_OUT), .A1 (N1451), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM415 (.ZN (XNOR_1_2_NAND2_NUM415_OUT), .A1 (GND), .A2 (N1492));
      NOR2_X1 XNOR_1_3_NAND2_NUM415 (.ZN (XNOR_1_3_NAND2_NUM415_OUT), .A1 (XNOR_1_1_NAND2_NUM415_OUT), .A2 (XNOR_1_2_NAND2_NUM415_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM415 (.ZN (N1520), .A1 (XNOR_1_3_NAND2_NUM415_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM416_OUT, XNOR_1_2_NAND2_NUM416_OUT, XNOR_1_3_NAND2_NUM416_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM416 (.ZN (XNOR_1_1_NAND2_NUM416_OUT), .A1 (N1453), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM416 (.ZN (XNOR_1_2_NAND2_NUM416_OUT), .A1 (GND), .A2 (N1493));
      NOR2_X1 XNOR_1_3_NAND2_NUM416 (.ZN (XNOR_1_3_NAND2_NUM416_OUT), .A1 (XNOR_1_1_NAND2_NUM416_OUT), .A2 (XNOR_1_2_NAND2_NUM416_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM416 (.ZN (N1521), .A1 (XNOR_1_3_NAND2_NUM416_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM417_OUT, XNOR_1_2_NAND2_NUM417_OUT, XNOR_1_3_NAND2_NUM417_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM417 (.ZN (XNOR_1_1_NAND2_NUM417_OUT), .A1 (N1455), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM417 (.ZN (XNOR_1_2_NAND2_NUM417_OUT), .A1 (GND), .A2 (N1494));
      NOR2_X1 XNOR_1_3_NAND2_NUM417 (.ZN (XNOR_1_3_NAND2_NUM417_OUT), .A1 (XNOR_1_1_NAND2_NUM417_OUT), .A2 (XNOR_1_2_NAND2_NUM417_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM417 (.ZN (N1522), .A1 (XNOR_1_3_NAND2_NUM417_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM418_OUT, XNOR_1_2_NAND2_NUM418_OUT, XNOR_1_3_NAND2_NUM418_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM418 (.ZN (XNOR_1_1_NAND2_NUM418_OUT), .A1 (N1457), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM418 (.ZN (XNOR_1_2_NAND2_NUM418_OUT), .A1 (GND), .A2 (N1495));
      NOR2_X1 XNOR_1_3_NAND2_NUM418 (.ZN (XNOR_1_3_NAND2_NUM418_OUT), .A1 (XNOR_1_1_NAND2_NUM418_OUT), .A2 (XNOR_1_2_NAND2_NUM418_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM418 (.ZN (N1526), .A1 (XNOR_1_3_NAND2_NUM418_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM419_OUT, XNOR_1_2_NAND2_NUM419_OUT, XNOR_1_3_NAND2_NUM419_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM419 (.ZN (XNOR_1_1_NAND2_NUM419_OUT), .A1 (N1459), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM419 (.ZN (XNOR_1_2_NAND2_NUM419_OUT), .A1 (GND), .A2 (N1496));
      NOR2_X1 XNOR_1_3_NAND2_NUM419 (.ZN (XNOR_1_3_NAND2_NUM419_OUT), .A1 (XNOR_1_1_NAND2_NUM419_OUT), .A2 (XNOR_1_2_NAND2_NUM419_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM419 (.ZN (N1527), .A1 (XNOR_1_3_NAND2_NUM419_OUT), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM420 (.ZN (N1528), .A1 (N1472), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM421_OUT, XNOR_1_2_NAND2_NUM421_OUT, XNOR_1_3_NAND2_NUM421_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM421 (.ZN (XNOR_1_1_NAND2_NUM421_OUT), .A1 (N1462), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM421 (.ZN (XNOR_1_2_NAND2_NUM421_OUT), .A1 (GND), .A2 (N1498));
      NOR2_X1 XNOR_1_3_NAND2_NUM421 (.ZN (XNOR_1_3_NAND2_NUM421_OUT), .A1 (XNOR_1_1_NAND2_NUM421_OUT), .A2 (XNOR_1_2_NAND2_NUM421_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM421 (.ZN (N1529), .A1 (XNOR_1_3_NAND2_NUM421_OUT), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM422 (.ZN (N1530), .A1 (N1478), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM423 (.ZN (N1531), .A1 (N1481), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM424 (.ZN (N1532), .A1 (N1484), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM425_OUT, XNOR_1_2_NAND2_NUM425_OUT, XNOR_1_3_NAND2_NUM425_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM425 (.ZN (XNOR_1_1_NAND2_NUM425_OUT), .A1 (N1471), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM425 (.ZN (XNOR_1_2_NAND2_NUM425_OUT), .A1 (GND), .A2 (N1501));
      NOR2_X1 XNOR_1_3_NAND2_NUM425 (.ZN (XNOR_1_3_NAND2_NUM425_OUT), .A1 (XNOR_1_1_NAND2_NUM425_OUT), .A2 (XNOR_1_2_NAND2_NUM425_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM425 (.ZN (N1534), .A1 (XNOR_1_3_NAND2_NUM425_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM426_OUT, XNOR_1_2_NAND2_NUM426_OUT, XNOR_1_3_NAND2_NUM426_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM426 (.ZN (XNOR_1_1_NAND2_NUM426_OUT), .A1 (N1469), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM426 (.ZN (XNOR_1_2_NAND2_NUM426_OUT), .A1 (GND), .A2 (N1500));
      NOR2_X1 XNOR_1_3_NAND2_NUM426 (.ZN (XNOR_1_3_NAND2_NUM426_OUT), .A1 (XNOR_1_1_NAND2_NUM426_OUT), .A2 (XNOR_1_2_NAND2_NUM426_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM426 (.ZN (N1537), .A1 (XNOR_1_3_NAND2_NUM426_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM427_OUT, XNOR_1_2_NAND2_NUM427_OUT, XNOR_1_3_NAND2_NUM427_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM427 (.ZN (XNOR_1_1_NAND2_NUM427_OUT), .A1 (N1476), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM427 (.ZN (XNOR_1_2_NAND2_NUM427_OUT), .A1 (GND), .A2 (N1504));
      NOR2_X1 XNOR_1_3_NAND2_NUM427 (.ZN (XNOR_1_3_NAND2_NUM427_OUT), .A1 (XNOR_1_1_NAND2_NUM427_OUT), .A2 (XNOR_1_2_NAND2_NUM427_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM427 (.ZN (N1540), .A1 (XNOR_1_3_NAND2_NUM427_OUT), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM428 (.ZN (N1546), .A1 (N1513), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM429 (.ZN (N1554), .A1 (N1521), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM430 (.ZN (N1557), .A1 (N1526), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM431 (.ZN (N1561), .A1 (N1520), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM432_OUT, XNOR_1_2_NAND2_NUM432_OUT, XNOR_1_3_NAND2_NUM432_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM432 (.ZN (XNOR_1_1_NAND2_NUM432_OUT), .A1 (N1484), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM432 (.ZN (XNOR_1_2_NAND2_NUM432_OUT), .A1 (GND), .A2 (N1531));
      NOR2_X1 XNOR_1_3_NAND2_NUM432 (.ZN (XNOR_1_3_NAND2_NUM432_OUT), .A1 (XNOR_1_1_NAND2_NUM432_OUT), .A2 (XNOR_1_2_NAND2_NUM432_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM432 (.ZN (N1567), .A1 (XNOR_1_3_NAND2_NUM432_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM433_OUT, XNOR_1_2_NAND2_NUM433_OUT, XNOR_1_3_NAND2_NUM433_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM433 (.ZN (XNOR_1_1_NAND2_NUM433_OUT), .A1 (N1481), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM433 (.ZN (XNOR_1_2_NAND2_NUM433_OUT), .A1 (GND), .A2 (N1532));
      NOR2_X1 XNOR_1_3_NAND2_NUM433 (.ZN (XNOR_1_3_NAND2_NUM433_OUT), .A1 (XNOR_1_1_NAND2_NUM433_OUT), .A2 (XNOR_1_2_NAND2_NUM433_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM433 (.ZN (N1568), .A1 (XNOR_1_3_NAND2_NUM433_OUT), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM434 (.ZN (N1569), .A1 (N1510), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM435 (.ZN (N1571), .A1 (N1527), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM436 (.ZN (N1576), .A1 (N1529), .A2 (GND));
      wire XNOR_1_1_BUFF1_NUM437_OUT;
      NOR2_X1 XNOR_1_1_BUFF1_NUM437 (.ZN (XNOR_1_1_BUFF1_NUM437_OUT), .A1 (N1522), .A2 (GND));
      NOR2_X1 XNOR_1_2_BUFF1_NUM437 (.ZN (N1588), .A1 (XNOR_1_1_BUFF1_NUM437_OUT), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM438 (.ZN (N1591), .A1 (N1534), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM439 (.ZN (N1593), .A1 (N1537), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM440_OUT, XNOR_1_2_NAND2_NUM440_OUT, XNOR_1_3_NAND2_NUM440_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM440 (.ZN (XNOR_1_1_NAND2_NUM440_OUT), .A1 (N1540), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM440 (.ZN (XNOR_1_2_NAND2_NUM440_OUT), .A1 (GND), .A2 (N1530));
      NOR2_X1 XNOR_1_3_NAND2_NUM440 (.ZN (XNOR_1_3_NAND2_NUM440_OUT), .A1 (XNOR_1_1_NAND2_NUM440_OUT), .A2 (XNOR_1_2_NAND2_NUM440_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM440 (.ZN (N1594), .A1 (XNOR_1_3_NAND2_NUM440_OUT), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM441 (.ZN (N1595), .A1 (N1540), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM442_OUT, XNOR_1_2_NAND2_NUM442_OUT, XNOR_1_3_NAND2_NUM442_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM442 (.ZN (XNOR_1_1_NAND2_NUM442_OUT), .A1 (N1567), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM442 (.ZN (XNOR_1_2_NAND2_NUM442_OUT), .A1 (GND), .A2 (N1568));
      NOR2_X1 XNOR_1_3_NAND2_NUM442 (.ZN (XNOR_1_3_NAND2_NUM442_OUT), .A1 (XNOR_1_1_NAND2_NUM442_OUT), .A2 (XNOR_1_2_NAND2_NUM442_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM442 (.ZN (N1596), .A1 (XNOR_1_3_NAND2_NUM442_OUT), .A2 (GND));
      wire XNOR_1_1_BUFF1_NUM443_OUT;
      NOR2_X1 XNOR_1_1_BUFF1_NUM443 (.ZN (XNOR_1_1_BUFF1_NUM443_OUT), .A1 (N1517), .A2 (GND));
      NOR2_X1 XNOR_1_2_BUFF1_NUM443 (.ZN (N1600), .A1 (XNOR_1_1_BUFF1_NUM443_OUT), .A2 (GND));
      wire XNOR_1_1_BUFF1_NUM444_OUT;
      NOR2_X1 XNOR_1_1_BUFF1_NUM444 (.ZN (XNOR_1_1_BUFF1_NUM444_OUT), .A1 (N1517), .A2 (GND));
      NOR2_X1 XNOR_1_2_BUFF1_NUM444 (.ZN (N1603), .A1 (XNOR_1_1_BUFF1_NUM444_OUT), .A2 (GND));
      wire XNOR_1_1_BUFF1_NUM445_OUT;
      NOR2_X1 XNOR_1_1_BUFF1_NUM445 (.ZN (XNOR_1_1_BUFF1_NUM445_OUT), .A1 (N1522), .A2 (GND));
      NOR2_X1 XNOR_1_2_BUFF1_NUM445 (.ZN (N1606), .A1 (XNOR_1_1_BUFF1_NUM445_OUT), .A2 (GND));
      wire XNOR_1_1_BUFF1_NUM446_OUT;
      NOR2_X1 XNOR_1_1_BUFF1_NUM446 (.ZN (XNOR_1_1_BUFF1_NUM446_OUT), .A1 (N1522), .A2 (GND));
      NOR2_X1 XNOR_1_2_BUFF1_NUM446 (.ZN (N1609), .A1 (XNOR_1_1_BUFF1_NUM446_OUT), .A2 (GND));
      wire XNOR_1_1_BUFF1_NUM447_OUT;
      NOR2_X1 XNOR_1_1_BUFF1_NUM447 (.ZN (XNOR_1_1_BUFF1_NUM447_OUT), .A1 (N1514), .A2 (GND));
      NOR2_X1 XNOR_1_2_BUFF1_NUM447 (.ZN (N1612), .A1 (XNOR_1_1_BUFF1_NUM447_OUT), .A2 (GND));
      wire XNOR_1_1_BUFF1_NUM448_OUT;
      NOR2_X1 XNOR_1_1_BUFF1_NUM448 (.ZN (XNOR_1_1_BUFF1_NUM448_OUT), .A1 (N1514), .A2 (GND));
      NOR2_X1 XNOR_1_2_BUFF1_NUM448 (.ZN (N1615), .A1 (XNOR_1_1_BUFF1_NUM448_OUT), .A2 (GND));
      wire XNOR_1_1_BUFF1_NUM449_OUT;
      NOR2_X1 XNOR_1_1_BUFF1_NUM449 (.ZN (XNOR_1_1_BUFF1_NUM449_OUT), .A1 (N1557), .A2 (GND));
      NOR2_X1 XNOR_1_2_BUFF1_NUM449 (.ZN (N1620), .A1 (XNOR_1_1_BUFF1_NUM449_OUT), .A2 (GND));
      wire XNOR_1_1_BUFF1_NUM450_OUT;
      NOR2_X1 XNOR_1_1_BUFF1_NUM450 (.ZN (XNOR_1_1_BUFF1_NUM450_OUT), .A1 (N1554), .A2 (GND));
      NOR2_X1 XNOR_1_2_BUFF1_NUM450 (.ZN (N1623), .A1 (XNOR_1_1_BUFF1_NUM450_OUT), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM451 (.ZN (N1635), .A1 (N1571), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM452_OUT, XNOR_1_2_NAND2_NUM452_OUT, XNOR_1_3_NAND2_NUM452_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM452 (.ZN (XNOR_1_1_NAND2_NUM452_OUT), .A1 (N1478), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM452 (.ZN (XNOR_1_2_NAND2_NUM452_OUT), .A1 (GND), .A2 (N1595));
      NOR2_X1 XNOR_1_3_NAND2_NUM452 (.ZN (XNOR_1_3_NAND2_NUM452_OUT), .A1 (XNOR_1_1_NAND2_NUM452_OUT), .A2 (XNOR_1_2_NAND2_NUM452_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM452 (.ZN (N1636), .A1 (XNOR_1_3_NAND2_NUM452_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM453_OUT, XNOR_1_2_NAND2_NUM453_OUT, XNOR_1_3_NAND2_NUM453_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM453 (.ZN (XNOR_1_1_NAND2_NUM453_OUT), .A1 (N1576), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM453 (.ZN (XNOR_1_2_NAND2_NUM453_OUT), .A1 (GND), .A2 (N1569));
      NOR2_X1 XNOR_1_3_NAND2_NUM453 (.ZN (XNOR_1_3_NAND2_NUM453_OUT), .A1 (XNOR_1_1_NAND2_NUM453_OUT), .A2 (XNOR_1_2_NAND2_NUM453_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM453 (.ZN (N1638), .A1 (XNOR_1_3_NAND2_NUM453_OUT), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM454 (.ZN (N1639), .A1 (N1576), .A2 (GND));
      wire XNOR_1_1_BUFF1_NUM455_OUT;
      NOR2_X1 XNOR_1_1_BUFF1_NUM455 (.ZN (XNOR_1_1_BUFF1_NUM455_OUT), .A1 (N1561), .A2 (GND));
      NOR2_X1 XNOR_1_2_BUFF1_NUM455 (.ZN (N1640), .A1 (XNOR_1_1_BUFF1_NUM455_OUT), .A2 (GND));
      wire XNOR_1_1_BUFF1_NUM456_OUT;
      NOR2_X1 XNOR_1_1_BUFF1_NUM456 (.ZN (XNOR_1_1_BUFF1_NUM456_OUT), .A1 (N1561), .A2 (GND));
      NOR2_X1 XNOR_1_2_BUFF1_NUM456 (.ZN (N1643), .A1 (XNOR_1_1_BUFF1_NUM456_OUT), .A2 (GND));
      wire XNOR_1_1_BUFF1_NUM457_OUT;
      NOR2_X1 XNOR_1_1_BUFF1_NUM457 (.ZN (XNOR_1_1_BUFF1_NUM457_OUT), .A1 (N1546), .A2 (GND));
      NOR2_X1 XNOR_1_2_BUFF1_NUM457 (.ZN (N1647), .A1 (XNOR_1_1_BUFF1_NUM457_OUT), .A2 (GND));
      wire XNOR_1_1_BUFF1_NUM458_OUT;
      NOR2_X1 XNOR_1_1_BUFF1_NUM458 (.ZN (XNOR_1_1_BUFF1_NUM458_OUT), .A1 (N1546), .A2 (GND));
      NOR2_X1 XNOR_1_2_BUFF1_NUM458 (.ZN (N1651), .A1 (XNOR_1_1_BUFF1_NUM458_OUT), .A2 (GND));
      wire XNOR_1_1_BUFF1_NUM459_OUT;
      NOR2_X1 XNOR_1_1_BUFF1_NUM459 (.ZN (XNOR_1_1_BUFF1_NUM459_OUT), .A1 (N1554), .A2 (GND));
      NOR2_X1 XNOR_1_2_BUFF1_NUM459 (.ZN (N1658), .A1 (XNOR_1_1_BUFF1_NUM459_OUT), .A2 (GND));
      wire XNOR_1_1_BUFF1_NUM460_OUT;
      NOR2_X1 XNOR_1_1_BUFF1_NUM460 (.ZN (XNOR_1_1_BUFF1_NUM460_OUT), .A1 (N1557), .A2 (GND));
      NOR2_X1 XNOR_1_2_BUFF1_NUM460 (.ZN (N1661), .A1 (XNOR_1_1_BUFF1_NUM460_OUT), .A2 (GND));
      wire XNOR_1_1_BUFF1_NUM461_OUT;
      NOR2_X1 XNOR_1_1_BUFF1_NUM461 (.ZN (XNOR_1_1_BUFF1_NUM461_OUT), .A1 (N1557), .A2 (GND));
      NOR2_X1 XNOR_1_2_BUFF1_NUM461 (.ZN (N1664), .A1 (XNOR_1_1_BUFF1_NUM461_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM462_OUT, XNOR_1_2_NAND2_NUM462_OUT, XNOR_1_3_NAND2_NUM462_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM462 (.ZN (XNOR_1_1_NAND2_NUM462_OUT), .A1 (N1596), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM462 (.ZN (XNOR_1_2_NAND2_NUM462_OUT), .A1 (GND), .A2 (N893));
      NOR2_X1 XNOR_1_3_NAND2_NUM462 (.ZN (XNOR_1_3_NAND2_NUM462_OUT), .A1 (XNOR_1_1_NAND2_NUM462_OUT), .A2 (XNOR_1_2_NAND2_NUM462_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM462 (.ZN (N1671), .A1 (XNOR_1_3_NAND2_NUM462_OUT), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM463 (.ZN (N1672), .A1 (N1596), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM464 (.ZN (N1675), .A1 (N1600), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM465 (.ZN (N1677), .A1 (N1603), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM466_OUT, XNOR_1_2_NAND2_NUM466_OUT, XNOR_1_3_NAND2_NUM466_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM466 (.ZN (XNOR_1_1_NAND2_NUM466_OUT), .A1 (N1606), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM466 (.ZN (XNOR_1_2_NAND2_NUM466_OUT), .A1 (GND), .A2 (N1217));
      NOR2_X1 XNOR_1_3_NAND2_NUM466 (.ZN (XNOR_1_3_NAND2_NUM466_OUT), .A1 (XNOR_1_1_NAND2_NUM466_OUT), .A2 (XNOR_1_2_NAND2_NUM466_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM466 (.ZN (N1678), .A1 (XNOR_1_3_NAND2_NUM466_OUT), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM467 (.ZN (N1679), .A1 (N1606), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM468_OUT, XNOR_1_2_NAND2_NUM468_OUT, XNOR_1_3_NAND2_NUM468_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM468 (.ZN (XNOR_1_1_NAND2_NUM468_OUT), .A1 (N1609), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM468 (.ZN (XNOR_1_2_NAND2_NUM468_OUT), .A1 (GND), .A2 (N1219));
      NOR2_X1 XNOR_1_3_NAND2_NUM468 (.ZN (XNOR_1_3_NAND2_NUM468_OUT), .A1 (XNOR_1_1_NAND2_NUM468_OUT), .A2 (XNOR_1_2_NAND2_NUM468_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM468 (.ZN (N1680), .A1 (XNOR_1_3_NAND2_NUM468_OUT), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM469 (.ZN (N1681), .A1 (N1609), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM470 (.ZN (N1682), .A1 (N1612), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM471 (.ZN (N1683), .A1 (N1615), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM472_OUT, XNOR_1_2_NAND2_NUM472_OUT, XNOR_1_3_NAND2_NUM472_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM472 (.ZN (XNOR_1_1_NAND2_NUM472_OUT), .A1 (N1594), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM472 (.ZN (XNOR_1_2_NAND2_NUM472_OUT), .A1 (GND), .A2 (N1636));
      NOR2_X1 XNOR_1_3_NAND2_NUM472 (.ZN (XNOR_1_3_NAND2_NUM472_OUT), .A1 (XNOR_1_1_NAND2_NUM472_OUT), .A2 (XNOR_1_2_NAND2_NUM472_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM472 (.ZN (N1685), .A1 (XNOR_1_3_NAND2_NUM472_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM473_OUT, XNOR_1_2_NAND2_NUM473_OUT, XNOR_1_3_NAND2_NUM473_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM473 (.ZN (XNOR_1_1_NAND2_NUM473_OUT), .A1 (N1510), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM473 (.ZN (XNOR_1_2_NAND2_NUM473_OUT), .A1 (GND), .A2 (N1639));
      NOR2_X1 XNOR_1_3_NAND2_NUM473 (.ZN (XNOR_1_3_NAND2_NUM473_OUT), .A1 (XNOR_1_1_NAND2_NUM473_OUT), .A2 (XNOR_1_2_NAND2_NUM473_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM473 (.ZN (N1688), .A1 (XNOR_1_3_NAND2_NUM473_OUT), .A2 (GND));
      wire XNOR_1_1_BUFF1_NUM474_OUT;
      NOR2_X1 XNOR_1_1_BUFF1_NUM474 (.ZN (XNOR_1_1_BUFF1_NUM474_OUT), .A1 (N1588), .A2 (GND));
      NOR2_X1 XNOR_1_2_BUFF1_NUM474 (.ZN (N1697), .A1 (XNOR_1_1_BUFF1_NUM474_OUT), .A2 (GND));
      wire XNOR_1_1_BUFF1_NUM475_OUT;
      NOR2_X1 XNOR_1_1_BUFF1_NUM475 (.ZN (XNOR_1_1_BUFF1_NUM475_OUT), .A1 (N1588), .A2 (GND));
      NOR2_X1 XNOR_1_2_BUFF1_NUM475 (.ZN (N1701), .A1 (XNOR_1_1_BUFF1_NUM475_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM476_OUT, XNOR_1_2_NAND2_NUM476_OUT, XNOR_1_3_NAND2_NUM476_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM476 (.ZN (XNOR_1_1_NAND2_NUM476_OUT), .A1 (N643), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM476 (.ZN (XNOR_1_2_NAND2_NUM476_OUT), .A1 (GND), .A2 (N1672));
      NOR2_X1 XNOR_1_3_NAND2_NUM476 (.ZN (XNOR_1_3_NAND2_NUM476_OUT), .A1 (XNOR_1_1_NAND2_NUM476_OUT), .A2 (XNOR_1_2_NAND2_NUM476_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM476 (.ZN (N1706), .A1 (XNOR_1_3_NAND2_NUM476_OUT), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM477 (.ZN (N1707), .A1 (N1643), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM478_OUT, XNOR_1_2_NAND2_NUM478_OUT, XNOR_1_3_NAND2_NUM478_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM478 (.ZN (XNOR_1_1_NAND2_NUM478_OUT), .A1 (N1647), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM478 (.ZN (XNOR_1_2_NAND2_NUM478_OUT), .A1 (GND), .A2 (N1675));
      NOR2_X1 XNOR_1_3_NAND2_NUM478 (.ZN (XNOR_1_3_NAND2_NUM478_OUT), .A1 (XNOR_1_1_NAND2_NUM478_OUT), .A2 (XNOR_1_2_NAND2_NUM478_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM478 (.ZN (N1708), .A1 (XNOR_1_3_NAND2_NUM478_OUT), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM479 (.ZN (N1709), .A1 (N1647), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM480_OUT, XNOR_1_2_NAND2_NUM480_OUT, XNOR_1_3_NAND2_NUM480_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM480 (.ZN (XNOR_1_1_NAND2_NUM480_OUT), .A1 (N1651), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM480 (.ZN (XNOR_1_2_NAND2_NUM480_OUT), .A1 (GND), .A2 (N1677));
      NOR2_X1 XNOR_1_3_NAND2_NUM480 (.ZN (XNOR_1_3_NAND2_NUM480_OUT), .A1 (XNOR_1_1_NAND2_NUM480_OUT), .A2 (XNOR_1_2_NAND2_NUM480_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM480 (.ZN (N1710), .A1 (XNOR_1_3_NAND2_NUM480_OUT), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM481 (.ZN (N1711), .A1 (N1651), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM482_OUT, XNOR_1_2_NAND2_NUM482_OUT, XNOR_1_3_NAND2_NUM482_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM482 (.ZN (XNOR_1_1_NAND2_NUM482_OUT), .A1 (N1028), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM482 (.ZN (XNOR_1_2_NAND2_NUM482_OUT), .A1 (GND), .A2 (N1679));
      NOR2_X1 XNOR_1_3_NAND2_NUM482 (.ZN (XNOR_1_3_NAND2_NUM482_OUT), .A1 (XNOR_1_1_NAND2_NUM482_OUT), .A2 (XNOR_1_2_NAND2_NUM482_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM482 (.ZN (N1712), .A1 (XNOR_1_3_NAND2_NUM482_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM483_OUT, XNOR_1_2_NAND2_NUM483_OUT, XNOR_1_3_NAND2_NUM483_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM483 (.ZN (XNOR_1_1_NAND2_NUM483_OUT), .A1 (N1031), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM483 (.ZN (XNOR_1_2_NAND2_NUM483_OUT), .A1 (GND), .A2 (N1681));
      NOR2_X1 XNOR_1_3_NAND2_NUM483 (.ZN (XNOR_1_3_NAND2_NUM483_OUT), .A1 (XNOR_1_1_NAND2_NUM483_OUT), .A2 (XNOR_1_2_NAND2_NUM483_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM483 (.ZN (N1713), .A1 (XNOR_1_3_NAND2_NUM483_OUT), .A2 (GND));
      wire XNOR_1_1_BUFF1_NUM484_OUT;
      NOR2_X1 XNOR_1_1_BUFF1_NUM484 (.ZN (XNOR_1_1_BUFF1_NUM484_OUT), .A1 (N1620), .A2 (GND));
      NOR2_X1 XNOR_1_2_BUFF1_NUM484 (.ZN (N1714), .A1 (XNOR_1_1_BUFF1_NUM484_OUT), .A2 (GND));
      wire XNOR_1_1_BUFF1_NUM485_OUT;
      NOR2_X1 XNOR_1_1_BUFF1_NUM485 (.ZN (XNOR_1_1_BUFF1_NUM485_OUT), .A1 (N1620), .A2 (GND));
      NOR2_X1 XNOR_1_2_BUFF1_NUM485 (.ZN (N1717), .A1 (XNOR_1_1_BUFF1_NUM485_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM486_OUT, XNOR_1_2_NAND2_NUM486_OUT, XNOR_1_3_NAND2_NUM486_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM486 (.ZN (XNOR_1_1_NAND2_NUM486_OUT), .A1 (N1658), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM486 (.ZN (XNOR_1_2_NAND2_NUM486_OUT), .A1 (GND), .A2 (N1593));
      NOR2_X1 XNOR_1_3_NAND2_NUM486 (.ZN (XNOR_1_3_NAND2_NUM486_OUT), .A1 (XNOR_1_1_NAND2_NUM486_OUT), .A2 (XNOR_1_2_NAND2_NUM486_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM486 (.ZN (N1720), .A1 (XNOR_1_3_NAND2_NUM486_OUT), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM487 (.ZN (N1721), .A1 (N1658), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM488_OUT, XNOR_1_2_NAND2_NUM488_OUT, XNOR_1_3_NAND2_NUM488_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM488 (.ZN (XNOR_1_1_NAND2_NUM488_OUT), .A1 (N1638), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM488 (.ZN (XNOR_1_2_NAND2_NUM488_OUT), .A1 (GND), .A2 (N1688));
      NOR2_X1 XNOR_1_3_NAND2_NUM488 (.ZN (XNOR_1_3_NAND2_NUM488_OUT), .A1 (XNOR_1_1_NAND2_NUM488_OUT), .A2 (XNOR_1_2_NAND2_NUM488_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM488 (.ZN (N1723), .A1 (XNOR_1_3_NAND2_NUM488_OUT), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM489 (.ZN (N1727), .A1 (N1661), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM490 (.ZN (N1728), .A1 (N1640), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM491 (.ZN (N1730), .A1 (N1664), .A2 (GND));
      wire XNOR_1_1_BUFF1_NUM492_OUT;
      NOR2_X1 XNOR_1_1_BUFF1_NUM492 (.ZN (XNOR_1_1_BUFF1_NUM492_OUT), .A1 (N1623), .A2 (GND));
      NOR2_X1 XNOR_1_2_BUFF1_NUM492 (.ZN (N1731), .A1 (XNOR_1_1_BUFF1_NUM492_OUT), .A2 (GND));
      wire XNOR_1_1_BUFF1_NUM493_OUT;
      NOR2_X1 XNOR_1_1_BUFF1_NUM493 (.ZN (XNOR_1_1_BUFF1_NUM493_OUT), .A1 (N1623), .A2 (GND));
      NOR2_X1 XNOR_1_2_BUFF1_NUM493 (.ZN (N1734), .A1 (XNOR_1_1_BUFF1_NUM493_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM494_OUT, XNOR_1_2_NAND2_NUM494_OUT, XNOR_1_3_NAND2_NUM494_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM494 (.ZN (XNOR_1_1_NAND2_NUM494_OUT), .A1 (N1685), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM494 (.ZN (XNOR_1_2_NAND2_NUM494_OUT), .A1 (GND), .A2 (N1528));
      NOR2_X1 XNOR_1_3_NAND2_NUM494 (.ZN (XNOR_1_3_NAND2_NUM494_OUT), .A1 (XNOR_1_1_NAND2_NUM494_OUT), .A2 (XNOR_1_2_NAND2_NUM494_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM494 (.ZN (N1740), .A1 (XNOR_1_3_NAND2_NUM494_OUT), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM495 (.ZN (N1741), .A1 (N1685), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM496_OUT, XNOR_1_2_NAND2_NUM496_OUT, XNOR_1_3_NAND2_NUM496_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM496 (.ZN (XNOR_1_1_NAND2_NUM496_OUT), .A1 (N1671), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM496 (.ZN (XNOR_1_2_NAND2_NUM496_OUT), .A1 (GND), .A2 (N1706));
      NOR2_X1 XNOR_1_3_NAND2_NUM496 (.ZN (XNOR_1_3_NAND2_NUM496_OUT), .A1 (XNOR_1_1_NAND2_NUM496_OUT), .A2 (XNOR_1_2_NAND2_NUM496_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM496 (.ZN (N1742), .A1 (XNOR_1_3_NAND2_NUM496_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM497_OUT, XNOR_1_2_NAND2_NUM497_OUT, XNOR_1_3_NAND2_NUM497_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM497 (.ZN (XNOR_1_1_NAND2_NUM497_OUT), .A1 (N1600), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM497 (.ZN (XNOR_1_2_NAND2_NUM497_OUT), .A1 (GND), .A2 (N1709));
      NOR2_X1 XNOR_1_3_NAND2_NUM497 (.ZN (XNOR_1_3_NAND2_NUM497_OUT), .A1 (XNOR_1_1_NAND2_NUM497_OUT), .A2 (XNOR_1_2_NAND2_NUM497_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM497 (.ZN (N1746), .A1 (XNOR_1_3_NAND2_NUM497_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM498_OUT, XNOR_1_2_NAND2_NUM498_OUT, XNOR_1_3_NAND2_NUM498_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM498 (.ZN (XNOR_1_1_NAND2_NUM498_OUT), .A1 (N1603), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM498 (.ZN (XNOR_1_2_NAND2_NUM498_OUT), .A1 (GND), .A2 (N1711));
      NOR2_X1 XNOR_1_3_NAND2_NUM498 (.ZN (XNOR_1_3_NAND2_NUM498_OUT), .A1 (XNOR_1_1_NAND2_NUM498_OUT), .A2 (XNOR_1_2_NAND2_NUM498_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM498 (.ZN (N1747), .A1 (XNOR_1_3_NAND2_NUM498_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM499_OUT, XNOR_1_2_NAND2_NUM499_OUT, XNOR_1_3_NAND2_NUM499_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM499 (.ZN (XNOR_1_1_NAND2_NUM499_OUT), .A1 (N1678), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM499 (.ZN (XNOR_1_2_NAND2_NUM499_OUT), .A1 (GND), .A2 (N1712));
      NOR2_X1 XNOR_1_3_NAND2_NUM499 (.ZN (XNOR_1_3_NAND2_NUM499_OUT), .A1 (XNOR_1_1_NAND2_NUM499_OUT), .A2 (XNOR_1_2_NAND2_NUM499_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM499 (.ZN (N1748), .A1 (XNOR_1_3_NAND2_NUM499_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM500_OUT, XNOR_1_2_NAND2_NUM500_OUT, XNOR_1_3_NAND2_NUM500_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM500 (.ZN (XNOR_1_1_NAND2_NUM500_OUT), .A1 (N1680), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM500 (.ZN (XNOR_1_2_NAND2_NUM500_OUT), .A1 (GND), .A2 (N1713));
      NOR2_X1 XNOR_1_3_NAND2_NUM500 (.ZN (XNOR_1_3_NAND2_NUM500_OUT), .A1 (XNOR_1_1_NAND2_NUM500_OUT), .A2 (XNOR_1_2_NAND2_NUM500_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM500 (.ZN (N1751), .A1 (XNOR_1_3_NAND2_NUM500_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM501_OUT, XNOR_1_2_NAND2_NUM501_OUT, XNOR_1_3_NAND2_NUM501_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM501 (.ZN (XNOR_1_1_NAND2_NUM501_OUT), .A1 (N1537), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM501 (.ZN (XNOR_1_2_NAND2_NUM501_OUT), .A1 (GND), .A2 (N1721));
      NOR2_X1 XNOR_1_3_NAND2_NUM501 (.ZN (XNOR_1_3_NAND2_NUM501_OUT), .A1 (XNOR_1_1_NAND2_NUM501_OUT), .A2 (XNOR_1_2_NAND2_NUM501_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM501 (.ZN (N1759), .A1 (XNOR_1_3_NAND2_NUM501_OUT), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM502 (.ZN (N1761), .A1 (N1697), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM503_OUT, XNOR_1_2_NAND2_NUM503_OUT, XNOR_1_3_NAND2_NUM503_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM503 (.ZN (XNOR_1_1_NAND2_NUM503_OUT), .A1 (N1697), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM503 (.ZN (XNOR_1_2_NAND2_NUM503_OUT), .A1 (GND), .A2 (N1727));
      NOR2_X1 XNOR_1_3_NAND2_NUM503 (.ZN (XNOR_1_3_NAND2_NUM503_OUT), .A1 (XNOR_1_1_NAND2_NUM503_OUT), .A2 (XNOR_1_2_NAND2_NUM503_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM503 (.ZN (N1762), .A1 (XNOR_1_3_NAND2_NUM503_OUT), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM504 (.ZN (N1763), .A1 (N1701), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM505_OUT, XNOR_1_2_NAND2_NUM505_OUT, XNOR_1_3_NAND2_NUM505_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM505 (.ZN (XNOR_1_1_NAND2_NUM505_OUT), .A1 (N1701), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM505 (.ZN (XNOR_1_2_NAND2_NUM505_OUT), .A1 (GND), .A2 (N1730));
      NOR2_X1 XNOR_1_3_NAND2_NUM505 (.ZN (XNOR_1_3_NAND2_NUM505_OUT), .A1 (XNOR_1_1_NAND2_NUM505_OUT), .A2 (XNOR_1_2_NAND2_NUM505_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM505 (.ZN (N1764), .A1 (XNOR_1_3_NAND2_NUM505_OUT), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM506 (.ZN (N1768), .A1 (N1717), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM507_OUT, XNOR_1_2_NAND2_NUM507_OUT, XNOR_1_3_NAND2_NUM507_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM507 (.ZN (XNOR_1_1_NAND2_NUM507_OUT), .A1 (N1472), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM507 (.ZN (XNOR_1_2_NAND2_NUM507_OUT), .A1 (GND), .A2 (N1741));
      NOR2_X1 XNOR_1_3_NAND2_NUM507 (.ZN (XNOR_1_3_NAND2_NUM507_OUT), .A1 (XNOR_1_1_NAND2_NUM507_OUT), .A2 (XNOR_1_2_NAND2_NUM507_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM507 (.ZN (N1769), .A1 (XNOR_1_3_NAND2_NUM507_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM508_OUT, XNOR_1_2_NAND2_NUM508_OUT, XNOR_1_3_NAND2_NUM508_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM508 (.ZN (XNOR_1_1_NAND2_NUM508_OUT), .A1 (N1723), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM508 (.ZN (XNOR_1_2_NAND2_NUM508_OUT), .A1 (GND), .A2 (N1413));
      NOR2_X1 XNOR_1_3_NAND2_NUM508 (.ZN (XNOR_1_3_NAND2_NUM508_OUT), .A1 (XNOR_1_1_NAND2_NUM508_OUT), .A2 (XNOR_1_2_NAND2_NUM508_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM508 (.ZN (N1772), .A1 (XNOR_1_3_NAND2_NUM508_OUT), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM509 (.ZN (N1773), .A1 (N1723), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM510_OUT, XNOR_1_2_NAND2_NUM510_OUT, XNOR_1_3_NAND2_NUM510_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM510 (.ZN (XNOR_1_1_NAND2_NUM510_OUT), .A1 (N1708), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM510 (.ZN (XNOR_1_2_NAND2_NUM510_OUT), .A1 (GND), .A2 (N1746));
      NOR2_X1 XNOR_1_3_NAND2_NUM510 (.ZN (XNOR_1_3_NAND2_NUM510_OUT), .A1 (XNOR_1_1_NAND2_NUM510_OUT), .A2 (XNOR_1_2_NAND2_NUM510_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM510 (.ZN (N1774), .A1 (XNOR_1_3_NAND2_NUM510_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM511_OUT, XNOR_1_2_NAND2_NUM511_OUT, XNOR_1_3_NAND2_NUM511_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM511 (.ZN (XNOR_1_1_NAND2_NUM511_OUT), .A1 (N1710), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM511 (.ZN (XNOR_1_2_NAND2_NUM511_OUT), .A1 (GND), .A2 (N1747));
      NOR2_X1 XNOR_1_3_NAND2_NUM511 (.ZN (XNOR_1_3_NAND2_NUM511_OUT), .A1 (XNOR_1_1_NAND2_NUM511_OUT), .A2 (XNOR_1_2_NAND2_NUM511_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM511 (.ZN (N1777), .A1 (XNOR_1_3_NAND2_NUM511_OUT), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM512 (.ZN (N1783), .A1 (N1731), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM513_OUT, XNOR_1_2_NAND2_NUM513_OUT, XNOR_1_3_NAND2_NUM513_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM513 (.ZN (XNOR_1_1_NAND2_NUM513_OUT), .A1 (N1731), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM513 (.ZN (XNOR_1_2_NAND2_NUM513_OUT), .A1 (GND), .A2 (N1682));
      NOR2_X1 XNOR_1_3_NAND2_NUM513 (.ZN (XNOR_1_3_NAND2_NUM513_OUT), .A1 (XNOR_1_1_NAND2_NUM513_OUT), .A2 (XNOR_1_2_NAND2_NUM513_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM513 (.ZN (N1784), .A1 (XNOR_1_3_NAND2_NUM513_OUT), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM514 (.ZN (N1785), .A1 (N1714), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM515 (.ZN (N1786), .A1 (N1734), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM516_OUT, XNOR_1_2_NAND2_NUM516_OUT, XNOR_1_3_NAND2_NUM516_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM516 (.ZN (XNOR_1_1_NAND2_NUM516_OUT), .A1 (N1734), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM516 (.ZN (XNOR_1_2_NAND2_NUM516_OUT), .A1 (GND), .A2 (N1683));
      NOR2_X1 XNOR_1_3_NAND2_NUM516 (.ZN (XNOR_1_3_NAND2_NUM516_OUT), .A1 (XNOR_1_1_NAND2_NUM516_OUT), .A2 (XNOR_1_2_NAND2_NUM516_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM516 (.ZN (N1787), .A1 (XNOR_1_3_NAND2_NUM516_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM517_OUT, XNOR_1_2_NAND2_NUM517_OUT, XNOR_1_3_NAND2_NUM517_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM517 (.ZN (XNOR_1_1_NAND2_NUM517_OUT), .A1 (N1720), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM517 (.ZN (XNOR_1_2_NAND2_NUM517_OUT), .A1 (GND), .A2 (N1759));
      NOR2_X1 XNOR_1_3_NAND2_NUM517 (.ZN (XNOR_1_3_NAND2_NUM517_OUT), .A1 (XNOR_1_1_NAND2_NUM517_OUT), .A2 (XNOR_1_2_NAND2_NUM517_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM517 (.ZN (N1788), .A1 (XNOR_1_3_NAND2_NUM517_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM518_OUT, XNOR_1_2_NAND2_NUM518_OUT, XNOR_1_3_NAND2_NUM518_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM518 (.ZN (XNOR_1_1_NAND2_NUM518_OUT), .A1 (N1661), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM518 (.ZN (XNOR_1_2_NAND2_NUM518_OUT), .A1 (GND), .A2 (N1761));
      NOR2_X1 XNOR_1_3_NAND2_NUM518 (.ZN (XNOR_1_3_NAND2_NUM518_OUT), .A1 (XNOR_1_1_NAND2_NUM518_OUT), .A2 (XNOR_1_2_NAND2_NUM518_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM518 (.ZN (N1791), .A1 (XNOR_1_3_NAND2_NUM518_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM519_OUT, XNOR_1_2_NAND2_NUM519_OUT, XNOR_1_3_NAND2_NUM519_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM519 (.ZN (XNOR_1_1_NAND2_NUM519_OUT), .A1 (N1664), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM519 (.ZN (XNOR_1_2_NAND2_NUM519_OUT), .A1 (GND), .A2 (N1763));
      NOR2_X1 XNOR_1_3_NAND2_NUM519 (.ZN (XNOR_1_3_NAND2_NUM519_OUT), .A1 (XNOR_1_1_NAND2_NUM519_OUT), .A2 (XNOR_1_2_NAND2_NUM519_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM519 (.ZN (N1792), .A1 (XNOR_1_3_NAND2_NUM519_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM520_OUT, XNOR_1_2_NAND2_NUM520_OUT, XNOR_1_3_NAND2_NUM520_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM520 (.ZN (XNOR_1_1_NAND2_NUM520_OUT), .A1 (N1751), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM520 (.ZN (XNOR_1_2_NAND2_NUM520_OUT), .A1 (GND), .A2 (N1155));
      NOR2_X1 XNOR_1_3_NAND2_NUM520 (.ZN (XNOR_1_3_NAND2_NUM520_OUT), .A1 (XNOR_1_1_NAND2_NUM520_OUT), .A2 (XNOR_1_2_NAND2_NUM520_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM520 (.ZN (N1795), .A1 (XNOR_1_3_NAND2_NUM520_OUT), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM521 (.ZN (N1796), .A1 (N1751), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM522_OUT, XNOR_1_2_NAND2_NUM522_OUT, XNOR_1_3_NAND2_NUM522_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM522 (.ZN (XNOR_1_1_NAND2_NUM522_OUT), .A1 (N1740), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM522 (.ZN (XNOR_1_2_NAND2_NUM522_OUT), .A1 (GND), .A2 (N1769));
      NOR2_X1 XNOR_1_3_NAND2_NUM522 (.ZN (XNOR_1_3_NAND2_NUM522_OUT), .A1 (XNOR_1_1_NAND2_NUM522_OUT), .A2 (XNOR_1_2_NAND2_NUM522_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM522 (.ZN (N1798), .A1 (XNOR_1_3_NAND2_NUM522_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM523_OUT, XNOR_1_2_NAND2_NUM523_OUT, XNOR_1_3_NAND2_NUM523_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM523 (.ZN (XNOR_1_1_NAND2_NUM523_OUT), .A1 (N1334), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM523 (.ZN (XNOR_1_2_NAND2_NUM523_OUT), .A1 (GND), .A2 (N1773));
      NOR2_X1 XNOR_1_3_NAND2_NUM523 (.ZN (XNOR_1_3_NAND2_NUM523_OUT), .A1 (XNOR_1_1_NAND2_NUM523_OUT), .A2 (XNOR_1_2_NAND2_NUM523_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM523 (.ZN (N1801), .A1 (XNOR_1_3_NAND2_NUM523_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM524_OUT, XNOR_1_2_NAND2_NUM524_OUT, XNOR_1_3_NAND2_NUM524_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM524 (.ZN (XNOR_1_1_NAND2_NUM524_OUT), .A1 (N1742), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM524 (.ZN (XNOR_1_2_NAND2_NUM524_OUT), .A1 (GND), .A2 (N290));
      NOR2_X1 XNOR_1_3_NAND2_NUM524 (.ZN (XNOR_1_3_NAND2_NUM524_OUT), .A1 (XNOR_1_1_NAND2_NUM524_OUT), .A2 (XNOR_1_2_NAND2_NUM524_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM524 (.ZN (N1802), .A1 (XNOR_1_3_NAND2_NUM524_OUT), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM525 (.ZN (N1807), .A1 (N1748), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM526_OUT, XNOR_1_2_NAND2_NUM526_OUT, XNOR_1_3_NAND2_NUM526_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM526 (.ZN (XNOR_1_1_NAND2_NUM526_OUT), .A1 (N1748), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM526 (.ZN (XNOR_1_2_NAND2_NUM526_OUT), .A1 (GND), .A2 (N1218));
      NOR2_X1 XNOR_1_3_NAND2_NUM526 (.ZN (XNOR_1_3_NAND2_NUM526_OUT), .A1 (XNOR_1_1_NAND2_NUM526_OUT), .A2 (XNOR_1_2_NAND2_NUM526_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM526 (.ZN (N1808), .A1 (XNOR_1_3_NAND2_NUM526_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM527_OUT, XNOR_1_2_NAND2_NUM527_OUT, XNOR_1_3_NAND2_NUM527_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM527 (.ZN (XNOR_1_1_NAND2_NUM527_OUT), .A1 (N1612), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM527 (.ZN (XNOR_1_2_NAND2_NUM527_OUT), .A1 (GND), .A2 (N1783));
      NOR2_X1 XNOR_1_3_NAND2_NUM527 (.ZN (XNOR_1_3_NAND2_NUM527_OUT), .A1 (XNOR_1_1_NAND2_NUM527_OUT), .A2 (XNOR_1_2_NAND2_NUM527_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM527 (.ZN (N1809), .A1 (XNOR_1_3_NAND2_NUM527_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM528_OUT, XNOR_1_2_NAND2_NUM528_OUT, XNOR_1_3_NAND2_NUM528_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM528 (.ZN (XNOR_1_1_NAND2_NUM528_OUT), .A1 (N1615), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM528 (.ZN (XNOR_1_2_NAND2_NUM528_OUT), .A1 (GND), .A2 (N1786));
      NOR2_X1 XNOR_1_3_NAND2_NUM528 (.ZN (XNOR_1_3_NAND2_NUM528_OUT), .A1 (XNOR_1_1_NAND2_NUM528_OUT), .A2 (XNOR_1_2_NAND2_NUM528_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM528 (.ZN (N1810), .A1 (XNOR_1_3_NAND2_NUM528_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM529_OUT, XNOR_1_2_NAND2_NUM529_OUT, XNOR_1_3_NAND2_NUM529_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM529 (.ZN (XNOR_1_1_NAND2_NUM529_OUT), .A1 (N1791), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM529 (.ZN (XNOR_1_2_NAND2_NUM529_OUT), .A1 (GND), .A2 (N1762));
      NOR2_X1 XNOR_1_3_NAND2_NUM529 (.ZN (XNOR_1_3_NAND2_NUM529_OUT), .A1 (XNOR_1_1_NAND2_NUM529_OUT), .A2 (XNOR_1_2_NAND2_NUM529_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM529 (.ZN (N1812), .A1 (XNOR_1_3_NAND2_NUM529_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM530_OUT, XNOR_1_2_NAND2_NUM530_OUT, XNOR_1_3_NAND2_NUM530_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM530 (.ZN (XNOR_1_1_NAND2_NUM530_OUT), .A1 (N1792), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM530 (.ZN (XNOR_1_2_NAND2_NUM530_OUT), .A1 (GND), .A2 (N1764));
      NOR2_X1 XNOR_1_3_NAND2_NUM530 (.ZN (XNOR_1_3_NAND2_NUM530_OUT), .A1 (XNOR_1_1_NAND2_NUM530_OUT), .A2 (XNOR_1_2_NAND2_NUM530_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM530 (.ZN (N1815), .A1 (XNOR_1_3_NAND2_NUM530_OUT), .A2 (GND));
      wire XNOR_1_1_BUFF1_NUM531_OUT;
      NOR2_X1 XNOR_1_1_BUFF1_NUM531 (.ZN (XNOR_1_1_BUFF1_NUM531_OUT), .A1 (N1742), .A2 (GND));
      NOR2_X1 XNOR_1_2_BUFF1_NUM531 (.ZN (N1818), .A1 (XNOR_1_1_BUFF1_NUM531_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM532_OUT, XNOR_1_2_NAND2_NUM532_OUT, XNOR_1_3_NAND2_NUM532_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM532 (.ZN (XNOR_1_1_NAND2_NUM532_OUT), .A1 (N1777), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM532 (.ZN (XNOR_1_2_NAND2_NUM532_OUT), .A1 (GND), .A2 (N1490));
      NOR2_X1 XNOR_1_3_NAND2_NUM532 (.ZN (XNOR_1_3_NAND2_NUM532_OUT), .A1 (XNOR_1_1_NAND2_NUM532_OUT), .A2 (XNOR_1_2_NAND2_NUM532_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM532 (.ZN (N1821), .A1 (XNOR_1_3_NAND2_NUM532_OUT), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM533 (.ZN (N1822), .A1 (N1777), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM534_OUT, XNOR_1_2_NAND2_NUM534_OUT, XNOR_1_3_NAND2_NUM534_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM534 (.ZN (XNOR_1_1_NAND2_NUM534_OUT), .A1 (N1774), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM534 (.ZN (XNOR_1_2_NAND2_NUM534_OUT), .A1 (GND), .A2 (N1491));
      NOR2_X1 XNOR_1_3_NAND2_NUM534 (.ZN (XNOR_1_3_NAND2_NUM534_OUT), .A1 (XNOR_1_1_NAND2_NUM534_OUT), .A2 (XNOR_1_2_NAND2_NUM534_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM534 (.ZN (N1823), .A1 (XNOR_1_3_NAND2_NUM534_OUT), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM535 (.ZN (N1824), .A1 (N1774), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM536_OUT, XNOR_1_2_NAND2_NUM536_OUT, XNOR_1_3_NAND2_NUM536_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM536 (.ZN (XNOR_1_1_NAND2_NUM536_OUT), .A1 (N962), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM536 (.ZN (XNOR_1_2_NAND2_NUM536_OUT), .A1 (GND), .A2 (N1796));
      NOR2_X1 XNOR_1_3_NAND2_NUM536 (.ZN (XNOR_1_3_NAND2_NUM536_OUT), .A1 (XNOR_1_1_NAND2_NUM536_OUT), .A2 (XNOR_1_2_NAND2_NUM536_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM536 (.ZN (N1825), .A1 (XNOR_1_3_NAND2_NUM536_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM537_OUT, XNOR_1_2_NAND2_NUM537_OUT, XNOR_1_3_NAND2_NUM537_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM537 (.ZN (XNOR_1_1_NAND2_NUM537_OUT), .A1 (N1788), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM537 (.ZN (XNOR_1_2_NAND2_NUM537_OUT), .A1 (GND), .A2 (N1409));
      NOR2_X1 XNOR_1_3_NAND2_NUM537 (.ZN (XNOR_1_3_NAND2_NUM537_OUT), .A1 (XNOR_1_1_NAND2_NUM537_OUT), .A2 (XNOR_1_2_NAND2_NUM537_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM537 (.ZN (N1826), .A1 (XNOR_1_3_NAND2_NUM537_OUT), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM538 (.ZN (N1827), .A1 (N1788), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM539_OUT, XNOR_1_2_NAND2_NUM539_OUT, XNOR_1_3_NAND2_NUM539_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM539 (.ZN (XNOR_1_1_NAND2_NUM539_OUT), .A1 (N1772), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM539 (.ZN (XNOR_1_2_NAND2_NUM539_OUT), .A1 (GND), .A2 (N1801));
      NOR2_X1 XNOR_1_3_NAND2_NUM539 (.ZN (XNOR_1_3_NAND2_NUM539_OUT), .A1 (XNOR_1_1_NAND2_NUM539_OUT), .A2 (XNOR_1_2_NAND2_NUM539_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM539 (.ZN (N1830), .A1 (XNOR_1_3_NAND2_NUM539_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM540_OUT, XNOR_1_2_NAND2_NUM540_OUT, XNOR_1_3_NAND2_NUM540_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM540 (.ZN (XNOR_1_1_NAND2_NUM540_OUT), .A1 (N959), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM540 (.ZN (XNOR_1_2_NAND2_NUM540_OUT), .A1 (GND), .A2 (N1807));
      NOR2_X1 XNOR_1_3_NAND2_NUM540 (.ZN (XNOR_1_3_NAND2_NUM540_OUT), .A1 (XNOR_1_1_NAND2_NUM540_OUT), .A2 (XNOR_1_2_NAND2_NUM540_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM540 (.ZN (N1837), .A1 (XNOR_1_3_NAND2_NUM540_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM541_OUT, XNOR_1_2_NAND2_NUM541_OUT, XNOR_1_3_NAND2_NUM541_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM541 (.ZN (XNOR_1_1_NAND2_NUM541_OUT), .A1 (N1809), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM541 (.ZN (XNOR_1_2_NAND2_NUM541_OUT), .A1 (GND), .A2 (N1784));
      NOR2_X1 XNOR_1_3_NAND2_NUM541 (.ZN (XNOR_1_3_NAND2_NUM541_OUT), .A1 (XNOR_1_1_NAND2_NUM541_OUT), .A2 (XNOR_1_2_NAND2_NUM541_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM541 (.ZN (N1838), .A1 (XNOR_1_3_NAND2_NUM541_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM542_OUT, XNOR_1_2_NAND2_NUM542_OUT, XNOR_1_3_NAND2_NUM542_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM542 (.ZN (XNOR_1_1_NAND2_NUM542_OUT), .A1 (N1810), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM542 (.ZN (XNOR_1_2_NAND2_NUM542_OUT), .A1 (GND), .A2 (N1787));
      NOR2_X1 XNOR_1_3_NAND2_NUM542 (.ZN (XNOR_1_3_NAND2_NUM542_OUT), .A1 (XNOR_1_1_NAND2_NUM542_OUT), .A2 (XNOR_1_2_NAND2_NUM542_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM542 (.ZN (N1841), .A1 (XNOR_1_3_NAND2_NUM542_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM543_OUT, XNOR_1_2_NAND2_NUM543_OUT, XNOR_1_3_NAND2_NUM543_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM543 (.ZN (XNOR_1_1_NAND2_NUM543_OUT), .A1 (N1419), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM543 (.ZN (XNOR_1_2_NAND2_NUM543_OUT), .A1 (GND), .A2 (N1822));
      NOR2_X1 XNOR_1_3_NAND2_NUM543 (.ZN (XNOR_1_3_NAND2_NUM543_OUT), .A1 (XNOR_1_1_NAND2_NUM543_OUT), .A2 (XNOR_1_2_NAND2_NUM543_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM543 (.ZN (N1848), .A1 (XNOR_1_3_NAND2_NUM543_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM544_OUT, XNOR_1_2_NAND2_NUM544_OUT, XNOR_1_3_NAND2_NUM544_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM544 (.ZN (XNOR_1_1_NAND2_NUM544_OUT), .A1 (N1416), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM544 (.ZN (XNOR_1_2_NAND2_NUM544_OUT), .A1 (GND), .A2 (N1824));
      NOR2_X1 XNOR_1_3_NAND2_NUM544 (.ZN (XNOR_1_3_NAND2_NUM544_OUT), .A1 (XNOR_1_1_NAND2_NUM544_OUT), .A2 (XNOR_1_2_NAND2_NUM544_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM544 (.ZN (N1849), .A1 (XNOR_1_3_NAND2_NUM544_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM545_OUT, XNOR_1_2_NAND2_NUM545_OUT, XNOR_1_3_NAND2_NUM545_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM545 (.ZN (XNOR_1_1_NAND2_NUM545_OUT), .A1 (N1795), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM545 (.ZN (XNOR_1_2_NAND2_NUM545_OUT), .A1 (GND), .A2 (N1825));
      NOR2_X1 XNOR_1_3_NAND2_NUM545 (.ZN (XNOR_1_3_NAND2_NUM545_OUT), .A1 (XNOR_1_1_NAND2_NUM545_OUT), .A2 (XNOR_1_2_NAND2_NUM545_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM545 (.ZN (N1850), .A1 (XNOR_1_3_NAND2_NUM545_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM546_OUT, XNOR_1_2_NAND2_NUM546_OUT, XNOR_1_3_NAND2_NUM546_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM546 (.ZN (XNOR_1_1_NAND2_NUM546_OUT), .A1 (N1319), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM546 (.ZN (XNOR_1_2_NAND2_NUM546_OUT), .A1 (GND), .A2 (N1827));
      NOR2_X1 XNOR_1_3_NAND2_NUM546 (.ZN (XNOR_1_3_NAND2_NUM546_OUT), .A1 (XNOR_1_1_NAND2_NUM546_OUT), .A2 (XNOR_1_2_NAND2_NUM546_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM546 (.ZN (N1852), .A1 (XNOR_1_3_NAND2_NUM546_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM547_OUT, XNOR_1_2_NAND2_NUM547_OUT, XNOR_1_3_NAND2_NUM547_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM547 (.ZN (XNOR_1_1_NAND2_NUM547_OUT), .A1 (N1815), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM547 (.ZN (XNOR_1_2_NAND2_NUM547_OUT), .A1 (GND), .A2 (N1707));
      NOR2_X1 XNOR_1_3_NAND2_NUM547 (.ZN (XNOR_1_3_NAND2_NUM547_OUT), .A1 (XNOR_1_1_NAND2_NUM547_OUT), .A2 (XNOR_1_2_NAND2_NUM547_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM547 (.ZN (N1855), .A1 (XNOR_1_3_NAND2_NUM547_OUT), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM548 (.ZN (N1856), .A1 (N1815), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM549 (.ZN (N1857), .A1 (N1818), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM550_OUT, XNOR_1_2_NAND2_NUM550_OUT, XNOR_1_3_NAND2_NUM550_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM550 (.ZN (XNOR_1_1_NAND2_NUM550_OUT), .A1 (N1798), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM550 (.ZN (XNOR_1_2_NAND2_NUM550_OUT), .A1 (GND), .A2 (N290));
      NOR2_X1 XNOR_1_3_NAND2_NUM550 (.ZN (XNOR_1_3_NAND2_NUM550_OUT), .A1 (XNOR_1_1_NAND2_NUM550_OUT), .A2 (XNOR_1_2_NAND2_NUM550_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM550 (.ZN (N1858), .A1 (XNOR_1_3_NAND2_NUM550_OUT), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM551 (.ZN (N1864), .A1 (N1812), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM552_OUT, XNOR_1_2_NAND2_NUM552_OUT, XNOR_1_3_NAND2_NUM552_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM552 (.ZN (XNOR_1_1_NAND2_NUM552_OUT), .A1 (N1812), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM552 (.ZN (XNOR_1_2_NAND2_NUM552_OUT), .A1 (GND), .A2 (N1728));
      NOR2_X1 XNOR_1_3_NAND2_NUM552 (.ZN (XNOR_1_3_NAND2_NUM552_OUT), .A1 (XNOR_1_1_NAND2_NUM552_OUT), .A2 (XNOR_1_2_NAND2_NUM552_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM552 (.ZN (N1865), .A1 (XNOR_1_3_NAND2_NUM552_OUT), .A2 (GND));
      wire XNOR_1_1_BUFF1_NUM553_OUT;
      NOR2_X1 XNOR_1_1_BUFF1_NUM553 (.ZN (XNOR_1_1_BUFF1_NUM553_OUT), .A1 (N1798), .A2 (GND));
      NOR2_X1 XNOR_1_2_BUFF1_NUM553 (.ZN (N1866), .A1 (XNOR_1_1_BUFF1_NUM553_OUT), .A2 (GND));
      wire XNOR_1_1_BUFF1_NUM554_OUT;
      NOR2_X1 XNOR_1_1_BUFF1_NUM554 (.ZN (XNOR_1_1_BUFF1_NUM554_OUT), .A1 (N1802), .A2 (GND));
      NOR2_X1 XNOR_1_2_BUFF1_NUM554 (.ZN (N1869), .A1 (XNOR_1_1_BUFF1_NUM554_OUT), .A2 (GND));
      wire XNOR_1_1_BUFF1_NUM555_OUT;
      NOR2_X1 XNOR_1_1_BUFF1_NUM555 (.ZN (XNOR_1_1_BUFF1_NUM555_OUT), .A1 (N1802), .A2 (GND));
      NOR2_X1 XNOR_1_2_BUFF1_NUM555 (.ZN (N1872), .A1 (XNOR_1_1_BUFF1_NUM555_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM556_OUT, XNOR_1_2_NAND2_NUM556_OUT, XNOR_1_3_NAND2_NUM556_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM556 (.ZN (XNOR_1_1_NAND2_NUM556_OUT), .A1 (N1808), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM556 (.ZN (XNOR_1_2_NAND2_NUM556_OUT), .A1 (GND), .A2 (N1837));
      NOR2_X1 XNOR_1_3_NAND2_NUM556 (.ZN (XNOR_1_3_NAND2_NUM556_OUT), .A1 (XNOR_1_1_NAND2_NUM556_OUT), .A2 (XNOR_1_2_NAND2_NUM556_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM556 (.ZN (N1875), .A1 (XNOR_1_3_NAND2_NUM556_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM557_OUT, XNOR_1_2_NAND2_NUM557_OUT, XNOR_1_3_NAND2_NUM557_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM557 (.ZN (XNOR_1_1_NAND2_NUM557_OUT), .A1 (N1821), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM557 (.ZN (XNOR_1_2_NAND2_NUM557_OUT), .A1 (GND), .A2 (N1848));
      NOR2_X1 XNOR_1_3_NAND2_NUM557 (.ZN (XNOR_1_3_NAND2_NUM557_OUT), .A1 (XNOR_1_1_NAND2_NUM557_OUT), .A2 (XNOR_1_2_NAND2_NUM557_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM557 (.ZN (N1878), .A1 (XNOR_1_3_NAND2_NUM557_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM558_OUT, XNOR_1_2_NAND2_NUM558_OUT, XNOR_1_3_NAND2_NUM558_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM558 (.ZN (XNOR_1_1_NAND2_NUM558_OUT), .A1 (N1823), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM558 (.ZN (XNOR_1_2_NAND2_NUM558_OUT), .A1 (GND), .A2 (N1849));
      NOR2_X1 XNOR_1_3_NAND2_NUM558 (.ZN (XNOR_1_3_NAND2_NUM558_OUT), .A1 (XNOR_1_1_NAND2_NUM558_OUT), .A2 (XNOR_1_2_NAND2_NUM558_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM558 (.ZN (N1879), .A1 (XNOR_1_3_NAND2_NUM558_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM559_OUT, XNOR_1_2_NAND2_NUM559_OUT, XNOR_1_3_NAND2_NUM559_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM559 (.ZN (XNOR_1_1_NAND2_NUM559_OUT), .A1 (N1841), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM559 (.ZN (XNOR_1_2_NAND2_NUM559_OUT), .A1 (GND), .A2 (N1768));
      NOR2_X1 XNOR_1_3_NAND2_NUM559 (.ZN (XNOR_1_3_NAND2_NUM559_OUT), .A1 (XNOR_1_1_NAND2_NUM559_OUT), .A2 (XNOR_1_2_NAND2_NUM559_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM559 (.ZN (N1882), .A1 (XNOR_1_3_NAND2_NUM559_OUT), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM560 (.ZN (N1883), .A1 (N1841), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM561_OUT, XNOR_1_2_NAND2_NUM561_OUT, XNOR_1_3_NAND2_NUM561_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM561 (.ZN (XNOR_1_1_NAND2_NUM561_OUT), .A1 (N1826), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM561 (.ZN (XNOR_1_2_NAND2_NUM561_OUT), .A1 (GND), .A2 (N1852));
      NOR2_X1 XNOR_1_3_NAND2_NUM561 (.ZN (XNOR_1_3_NAND2_NUM561_OUT), .A1 (XNOR_1_1_NAND2_NUM561_OUT), .A2 (XNOR_1_2_NAND2_NUM561_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM561 (.ZN (N1884), .A1 (XNOR_1_3_NAND2_NUM561_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM562_OUT, XNOR_1_2_NAND2_NUM562_OUT, XNOR_1_3_NAND2_NUM562_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM562 (.ZN (XNOR_1_1_NAND2_NUM562_OUT), .A1 (N1643), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM562 (.ZN (XNOR_1_2_NAND2_NUM562_OUT), .A1 (GND), .A2 (N1856));
      NOR2_X1 XNOR_1_3_NAND2_NUM562 (.ZN (XNOR_1_3_NAND2_NUM562_OUT), .A1 (XNOR_1_1_NAND2_NUM562_OUT), .A2 (XNOR_1_2_NAND2_NUM562_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM562 (.ZN (N1885), .A1 (XNOR_1_3_NAND2_NUM562_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM563_OUT, XNOR_1_2_NAND2_NUM563_OUT, XNOR_1_3_NAND2_NUM563_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM563 (.ZN (XNOR_1_1_NAND2_NUM563_OUT), .A1 (N1830), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM563 (.ZN (XNOR_1_2_NAND2_NUM563_OUT), .A1 (GND), .A2 (N290));
      NOR2_X1 XNOR_1_3_NAND2_NUM563 (.ZN (XNOR_1_3_NAND2_NUM563_OUT), .A1 (XNOR_1_1_NAND2_NUM563_OUT), .A2 (XNOR_1_2_NAND2_NUM563_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM563 (.ZN (N1889), .A1 (XNOR_1_3_NAND2_NUM563_OUT), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM564 (.ZN (N1895), .A1 (N1838), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM565_OUT, XNOR_1_2_NAND2_NUM565_OUT, XNOR_1_3_NAND2_NUM565_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM565 (.ZN (XNOR_1_1_NAND2_NUM565_OUT), .A1 (N1838), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM565 (.ZN (XNOR_1_2_NAND2_NUM565_OUT), .A1 (GND), .A2 (N1785));
      NOR2_X1 XNOR_1_3_NAND2_NUM565 (.ZN (XNOR_1_3_NAND2_NUM565_OUT), .A1 (XNOR_1_1_NAND2_NUM565_OUT), .A2 (XNOR_1_2_NAND2_NUM565_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM565 (.ZN (N1896), .A1 (XNOR_1_3_NAND2_NUM565_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM566_OUT, XNOR_1_2_NAND2_NUM566_OUT, XNOR_1_3_NAND2_NUM566_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM566 (.ZN (XNOR_1_1_NAND2_NUM566_OUT), .A1 (N1640), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM566 (.ZN (XNOR_1_2_NAND2_NUM566_OUT), .A1 (GND), .A2 (N1864));
      NOR2_X1 XNOR_1_3_NAND2_NUM566 (.ZN (XNOR_1_3_NAND2_NUM566_OUT), .A1 (XNOR_1_1_NAND2_NUM566_OUT), .A2 (XNOR_1_2_NAND2_NUM566_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM566 (.ZN (N1897), .A1 (XNOR_1_3_NAND2_NUM566_OUT), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM567 (.ZN (N1898), .A1 (N1850), .A2 (GND));
      wire XNOR_1_1_BUFF1_NUM568_OUT;
      NOR2_X1 XNOR_1_1_BUFF1_NUM568 (.ZN (XNOR_1_1_BUFF1_NUM568_OUT), .A1 (N1830), .A2 (GND));
      NOR2_X1 XNOR_1_2_BUFF1_NUM568 (.ZN (N1902), .A1 (XNOR_1_1_BUFF1_NUM568_OUT), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM569 (.ZN (N1910), .A1 (N1878), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM570_OUT, XNOR_1_2_NAND2_NUM570_OUT, XNOR_1_3_NAND2_NUM570_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM570 (.ZN (XNOR_1_1_NAND2_NUM570_OUT), .A1 (N1717), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM570 (.ZN (XNOR_1_2_NAND2_NUM570_OUT), .A1 (GND), .A2 (N1883));
      NOR2_X1 XNOR_1_3_NAND2_NUM570 (.ZN (XNOR_1_3_NAND2_NUM570_OUT), .A1 (XNOR_1_1_NAND2_NUM570_OUT), .A2 (XNOR_1_2_NAND2_NUM570_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM570 (.ZN (N1911), .A1 (XNOR_1_3_NAND2_NUM570_OUT), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM571 (.ZN (N1912), .A1 (N1884), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM572_OUT, XNOR_1_2_NAND2_NUM572_OUT, XNOR_1_3_NAND2_NUM572_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM572 (.ZN (XNOR_1_1_NAND2_NUM572_OUT), .A1 (N1855), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM572 (.ZN (XNOR_1_2_NAND2_NUM572_OUT), .A1 (GND), .A2 (N1885));
      NOR2_X1 XNOR_1_3_NAND2_NUM572 (.ZN (XNOR_1_3_NAND2_NUM572_OUT), .A1 (XNOR_1_1_NAND2_NUM572_OUT), .A2 (XNOR_1_2_NAND2_NUM572_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM572 (.ZN (N1913), .A1 (XNOR_1_3_NAND2_NUM572_OUT), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM573 (.ZN (N1915), .A1 (N1866), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM574_OUT, XNOR_1_2_NAND2_NUM574_OUT, XNOR_1_3_NAND2_NUM574_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM574 (.ZN (XNOR_1_1_NAND2_NUM574_OUT), .A1 (N1872), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM574 (.ZN (XNOR_1_2_NAND2_NUM574_OUT), .A1 (GND), .A2 (N919));
      NOR2_X1 XNOR_1_3_NAND2_NUM574 (.ZN (XNOR_1_3_NAND2_NUM574_OUT), .A1 (XNOR_1_1_NAND2_NUM574_OUT), .A2 (XNOR_1_2_NAND2_NUM574_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM574 (.ZN (N1919), .A1 (XNOR_1_3_NAND2_NUM574_OUT), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM575 (.ZN (N1920), .A1 (N1872), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM576_OUT, XNOR_1_2_NAND2_NUM576_OUT, XNOR_1_3_NAND2_NUM576_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM576 (.ZN (XNOR_1_1_NAND2_NUM576_OUT), .A1 (N1869), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM576 (.ZN (XNOR_1_2_NAND2_NUM576_OUT), .A1 (GND), .A2 (N920));
      NOR2_X1 XNOR_1_3_NAND2_NUM576 (.ZN (XNOR_1_3_NAND2_NUM576_OUT), .A1 (XNOR_1_1_NAND2_NUM576_OUT), .A2 (XNOR_1_2_NAND2_NUM576_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM576 (.ZN (N1921), .A1 (XNOR_1_3_NAND2_NUM576_OUT), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM577 (.ZN (N1922), .A1 (N1869), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM578 (.ZN (N1923), .A1 (N1875), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM579_OUT, XNOR_1_2_NAND2_NUM579_OUT, XNOR_1_3_NAND2_NUM579_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM579 (.ZN (XNOR_1_1_NAND2_NUM579_OUT), .A1 (N1714), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM579 (.ZN (XNOR_1_2_NAND2_NUM579_OUT), .A1 (GND), .A2 (N1895));
      NOR2_X1 XNOR_1_3_NAND2_NUM579 (.ZN (XNOR_1_3_NAND2_NUM579_OUT), .A1 (XNOR_1_1_NAND2_NUM579_OUT), .A2 (XNOR_1_2_NAND2_NUM579_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM579 (.ZN (N1924), .A1 (XNOR_1_3_NAND2_NUM579_OUT), .A2 (GND));
      wire XNOR_1_1_BUFF1_NUM580_OUT;
      NOR2_X1 XNOR_1_1_BUFF1_NUM580 (.ZN (XNOR_1_1_BUFF1_NUM580_OUT), .A1 (N1858), .A2 (GND));
      NOR2_X1 XNOR_1_2_BUFF1_NUM580 (.ZN (N1927), .A1 (XNOR_1_1_BUFF1_NUM580_OUT), .A2 (GND));
      wire XNOR_1_1_BUFF1_NUM581_OUT;
      NOR2_X1 XNOR_1_1_BUFF1_NUM581 (.ZN (XNOR_1_1_BUFF1_NUM581_OUT), .A1 (N1858), .A2 (GND));
      NOR2_X1 XNOR_1_2_BUFF1_NUM581 (.ZN (N1930), .A1 (XNOR_1_1_BUFF1_NUM581_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM582_OUT, XNOR_1_2_NAND2_NUM582_OUT, XNOR_1_3_NAND2_NUM582_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM582 (.ZN (XNOR_1_1_NAND2_NUM582_OUT), .A1 (N1865), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM582 (.ZN (XNOR_1_2_NAND2_NUM582_OUT), .A1 (GND), .A2 (N1897));
      NOR2_X1 XNOR_1_3_NAND2_NUM582 (.ZN (XNOR_1_3_NAND2_NUM582_OUT), .A1 (XNOR_1_1_NAND2_NUM582_OUT), .A2 (XNOR_1_2_NAND2_NUM582_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM582 (.ZN (N1933), .A1 (XNOR_1_3_NAND2_NUM582_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM583_OUT, XNOR_1_2_NAND2_NUM583_OUT, XNOR_1_3_NAND2_NUM583_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM583 (.ZN (XNOR_1_1_NAND2_NUM583_OUT), .A1 (N1882), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM583 (.ZN (XNOR_1_2_NAND2_NUM583_OUT), .A1 (GND), .A2 (N1911));
      NOR2_X1 XNOR_1_3_NAND2_NUM583 (.ZN (XNOR_1_3_NAND2_NUM583_OUT), .A1 (XNOR_1_1_NAND2_NUM583_OUT), .A2 (XNOR_1_2_NAND2_NUM583_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM583 (.ZN (N1936), .A1 (XNOR_1_3_NAND2_NUM583_OUT), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM584 (.ZN (N1937), .A1 (N1898), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM585 (.ZN (N1938), .A1 (N1902), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM586_OUT, XNOR_1_2_NAND2_NUM586_OUT, XNOR_1_3_NAND2_NUM586_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM586 (.ZN (XNOR_1_1_NAND2_NUM586_OUT), .A1 (N679), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM586 (.ZN (XNOR_1_2_NAND2_NUM586_OUT), .A1 (GND), .A2 (N1920));
      NOR2_X1 XNOR_1_3_NAND2_NUM586 (.ZN (XNOR_1_3_NAND2_NUM586_OUT), .A1 (XNOR_1_1_NAND2_NUM586_OUT), .A2 (XNOR_1_2_NAND2_NUM586_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM586 (.ZN (N1941), .A1 (XNOR_1_3_NAND2_NUM586_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM587_OUT, XNOR_1_2_NAND2_NUM587_OUT, XNOR_1_3_NAND2_NUM587_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM587 (.ZN (XNOR_1_1_NAND2_NUM587_OUT), .A1 (N676), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM587 (.ZN (XNOR_1_2_NAND2_NUM587_OUT), .A1 (GND), .A2 (N1922));
      NOR2_X1 XNOR_1_3_NAND2_NUM587 (.ZN (XNOR_1_3_NAND2_NUM587_OUT), .A1 (XNOR_1_1_NAND2_NUM587_OUT), .A2 (XNOR_1_2_NAND2_NUM587_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM587 (.ZN (N1942), .A1 (XNOR_1_3_NAND2_NUM587_OUT), .A2 (GND));
      wire XNOR_1_1_BUFF1_NUM588_OUT;
      NOR2_X1 XNOR_1_1_BUFF1_NUM588 (.ZN (XNOR_1_1_BUFF1_NUM588_OUT), .A1 (N1879), .A2 (GND));
      NOR2_X1 XNOR_1_2_BUFF1_NUM588 (.ZN (N1944), .A1 (XNOR_1_1_BUFF1_NUM588_OUT), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM589 (.ZN (N1947), .A1 (N1913), .A2 (GND));
      wire XNOR_1_1_BUFF1_NUM590_OUT;
      NOR2_X1 XNOR_1_1_BUFF1_NUM590 (.ZN (XNOR_1_1_BUFF1_NUM590_OUT), .A1 (N1889), .A2 (GND));
      NOR2_X1 XNOR_1_2_BUFF1_NUM590 (.ZN (N1950), .A1 (XNOR_1_1_BUFF1_NUM590_OUT), .A2 (GND));
      wire XNOR_1_1_BUFF1_NUM591_OUT;
      NOR2_X1 XNOR_1_1_BUFF1_NUM591 (.ZN (XNOR_1_1_BUFF1_NUM591_OUT), .A1 (N1889), .A2 (GND));
      NOR2_X1 XNOR_1_2_BUFF1_NUM591 (.ZN (N1953), .A1 (XNOR_1_1_BUFF1_NUM591_OUT), .A2 (GND));
      wire XNOR_1_1_BUFF1_NUM592_OUT;
      NOR2_X1 XNOR_1_1_BUFF1_NUM592 (.ZN (XNOR_1_1_BUFF1_NUM592_OUT), .A1 (N1879), .A2 (GND));
      NOR2_X1 XNOR_1_2_BUFF1_NUM592 (.ZN (N1958), .A1 (XNOR_1_1_BUFF1_NUM592_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM593_OUT, XNOR_1_2_NAND2_NUM593_OUT, XNOR_1_3_NAND2_NUM593_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM593 (.ZN (XNOR_1_1_NAND2_NUM593_OUT), .A1 (N1896), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM593 (.ZN (XNOR_1_2_NAND2_NUM593_OUT), .A1 (GND), .A2 (N1924));
      NOR2_X1 XNOR_1_3_NAND2_NUM593 (.ZN (XNOR_1_3_NAND2_NUM593_OUT), .A1 (XNOR_1_1_NAND2_NUM593_OUT), .A2 (XNOR_1_2_NAND2_NUM593_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM593 (.ZN (N1961), .A1 (XNOR_1_3_NAND2_NUM593_OUT), .A2 (GND));
      wire XNOR_1_1_AND2_NUM594_OUT, XNOR_1_2_AND2_NUM594_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM594 (.ZN (XNOR_1_1_AND2_NUM594_OUT), .A1 (N1910), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM594 (.ZN (XNOR_1_2_AND2_NUM594_OUT), .A1 (GND), .A2 (N601));
      NOR2_X1 XNOR_1_3_AND2_NUM594 (.ZN (N1965), .A1 (XNOR_1_1_AND2_NUM594_OUT), .A2 (XNOR_1_2_AND2_NUM594_OUT));
      wire XNOR_1_1_AND2_NUM595_OUT, XNOR_1_2_AND2_NUM595_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM595 (.ZN (XNOR_1_1_AND2_NUM595_OUT), .A1 (N602), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM595 (.ZN (XNOR_1_2_AND2_NUM595_OUT), .A1 (GND), .A2 (N1912));
      NOR2_X1 XNOR_1_3_AND2_NUM595 (.ZN (N1968), .A1 (XNOR_1_1_AND2_NUM595_OUT), .A2 (XNOR_1_2_AND2_NUM595_OUT));
      wire XNOR_1_1_NAND2_NUM596_OUT, XNOR_1_2_NAND2_NUM596_OUT, XNOR_1_3_NAND2_NUM596_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM596 (.ZN (XNOR_1_1_NAND2_NUM596_OUT), .A1 (N1930), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM596 (.ZN (XNOR_1_2_NAND2_NUM596_OUT), .A1 (GND), .A2 (N917));
      NOR2_X1 XNOR_1_3_NAND2_NUM596 (.ZN (XNOR_1_3_NAND2_NUM596_OUT), .A1 (XNOR_1_1_NAND2_NUM596_OUT), .A2 (XNOR_1_2_NAND2_NUM596_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM596 (.ZN (N1975), .A1 (XNOR_1_3_NAND2_NUM596_OUT), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM597 (.ZN (N1976), .A1 (N1930), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM598_OUT, XNOR_1_2_NAND2_NUM598_OUT, XNOR_1_3_NAND2_NUM598_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM598 (.ZN (XNOR_1_1_NAND2_NUM598_OUT), .A1 (N1927), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM598 (.ZN (XNOR_1_2_NAND2_NUM598_OUT), .A1 (GND), .A2 (N918));
      NOR2_X1 XNOR_1_3_NAND2_NUM598 (.ZN (XNOR_1_3_NAND2_NUM598_OUT), .A1 (XNOR_1_1_NAND2_NUM598_OUT), .A2 (XNOR_1_2_NAND2_NUM598_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM598 (.ZN (N1977), .A1 (XNOR_1_3_NAND2_NUM598_OUT), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM599 (.ZN (N1978), .A1 (N1927), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM600_OUT, XNOR_1_2_NAND2_NUM600_OUT, XNOR_1_3_NAND2_NUM600_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM600 (.ZN (XNOR_1_1_NAND2_NUM600_OUT), .A1 (N1919), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM600 (.ZN (XNOR_1_2_NAND2_NUM600_OUT), .A1 (GND), .A2 (N1941));
      NOR2_X1 XNOR_1_3_NAND2_NUM600 (.ZN (XNOR_1_3_NAND2_NUM600_OUT), .A1 (XNOR_1_1_NAND2_NUM600_OUT), .A2 (XNOR_1_2_NAND2_NUM600_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM600 (.ZN (N1979), .A1 (XNOR_1_3_NAND2_NUM600_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM601_OUT, XNOR_1_2_NAND2_NUM601_OUT, XNOR_1_3_NAND2_NUM601_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM601 (.ZN (XNOR_1_1_NAND2_NUM601_OUT), .A1 (N1921), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM601 (.ZN (XNOR_1_2_NAND2_NUM601_OUT), .A1 (GND), .A2 (N1942));
      NOR2_X1 XNOR_1_3_NAND2_NUM601 (.ZN (XNOR_1_3_NAND2_NUM601_OUT), .A1 (XNOR_1_1_NAND2_NUM601_OUT), .A2 (XNOR_1_2_NAND2_NUM601_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM601 (.ZN (N1980), .A1 (XNOR_1_3_NAND2_NUM601_OUT), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM602 (.ZN (N1985), .A1 (N1933), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM603 (.ZN (N1987), .A1 (N1936), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM604 (.ZN (N1999), .A1 (N1944), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM605_OUT, XNOR_1_2_NAND2_NUM605_OUT, XNOR_1_3_NAND2_NUM605_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM605 (.ZN (XNOR_1_1_NAND2_NUM605_OUT), .A1 (N1944), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM605 (.ZN (XNOR_1_2_NAND2_NUM605_OUT), .A1 (GND), .A2 (N1937));
      NOR2_X1 XNOR_1_3_NAND2_NUM605 (.ZN (XNOR_1_3_NAND2_NUM605_OUT), .A1 (XNOR_1_1_NAND2_NUM605_OUT), .A2 (XNOR_1_2_NAND2_NUM605_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM605 (.ZN (N2000), .A1 (XNOR_1_3_NAND2_NUM605_OUT), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM606 (.ZN (N2002), .A1 (N1947), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM607_OUT, XNOR_1_2_NAND2_NUM607_OUT, XNOR_1_3_NAND2_NUM607_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM607 (.ZN (XNOR_1_1_NAND2_NUM607_OUT), .A1 (N1947), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM607 (.ZN (XNOR_1_2_NAND2_NUM607_OUT), .A1 (GND), .A2 (N1499));
      NOR2_X1 XNOR_1_3_NAND2_NUM607 (.ZN (XNOR_1_3_NAND2_NUM607_OUT), .A1 (XNOR_1_1_NAND2_NUM607_OUT), .A2 (XNOR_1_2_NAND2_NUM607_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM607 (.ZN (N2003), .A1 (XNOR_1_3_NAND2_NUM607_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM608_OUT, XNOR_1_2_NAND2_NUM608_OUT, XNOR_1_3_NAND2_NUM608_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM608 (.ZN (XNOR_1_1_NAND2_NUM608_OUT), .A1 (N1953), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM608 (.ZN (XNOR_1_2_NAND2_NUM608_OUT), .A1 (GND), .A2 (N1350));
      NOR2_X1 XNOR_1_3_NAND2_NUM608 (.ZN (XNOR_1_3_NAND2_NUM608_OUT), .A1 (XNOR_1_1_NAND2_NUM608_OUT), .A2 (XNOR_1_2_NAND2_NUM608_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM608 (.ZN (N2004), .A1 (XNOR_1_3_NAND2_NUM608_OUT), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM609 (.ZN (N2005), .A1 (N1953), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM610_OUT, XNOR_1_2_NAND2_NUM610_OUT, XNOR_1_3_NAND2_NUM610_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM610 (.ZN (XNOR_1_1_NAND2_NUM610_OUT), .A1 (N1950), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM610 (.ZN (XNOR_1_2_NAND2_NUM610_OUT), .A1 (GND), .A2 (N1351));
      NOR2_X1 XNOR_1_3_NAND2_NUM610 (.ZN (XNOR_1_3_NAND2_NUM610_OUT), .A1 (XNOR_1_1_NAND2_NUM610_OUT), .A2 (XNOR_1_2_NAND2_NUM610_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM610 (.ZN (N2006), .A1 (XNOR_1_3_NAND2_NUM610_OUT), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM611 (.ZN (N2007), .A1 (N1950), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM612_OUT, XNOR_1_2_NAND2_NUM612_OUT, XNOR_1_3_NAND2_NUM612_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM612 (.ZN (XNOR_1_1_NAND2_NUM612_OUT), .A1 (N673), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM612 (.ZN (XNOR_1_2_NAND2_NUM612_OUT), .A1 (GND), .A2 (N1976));
      NOR2_X1 XNOR_1_3_NAND2_NUM612 (.ZN (XNOR_1_3_NAND2_NUM612_OUT), .A1 (XNOR_1_1_NAND2_NUM612_OUT), .A2 (XNOR_1_2_NAND2_NUM612_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM612 (.ZN (N2008), .A1 (XNOR_1_3_NAND2_NUM612_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM613_OUT, XNOR_1_2_NAND2_NUM613_OUT, XNOR_1_3_NAND2_NUM613_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM613 (.ZN (XNOR_1_1_NAND2_NUM613_OUT), .A1 (N670), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM613 (.ZN (XNOR_1_2_NAND2_NUM613_OUT), .A1 (GND), .A2 (N1978));
      NOR2_X1 XNOR_1_3_NAND2_NUM613 (.ZN (XNOR_1_3_NAND2_NUM613_OUT), .A1 (XNOR_1_1_NAND2_NUM613_OUT), .A2 (XNOR_1_2_NAND2_NUM613_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM613 (.ZN (N2009), .A1 (XNOR_1_3_NAND2_NUM613_OUT), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM614 (.ZN (N2012), .A1 (N1979), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM615 (.ZN (N2013), .A1 (N1958), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM616_OUT, XNOR_1_2_NAND2_NUM616_OUT, XNOR_1_3_NAND2_NUM616_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM616 (.ZN (XNOR_1_1_NAND2_NUM616_OUT), .A1 (N1958), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM616 (.ZN (XNOR_1_2_NAND2_NUM616_OUT), .A1 (GND), .A2 (N1923));
      NOR2_X1 XNOR_1_3_NAND2_NUM616 (.ZN (XNOR_1_3_NAND2_NUM616_OUT), .A1 (XNOR_1_1_NAND2_NUM616_OUT), .A2 (XNOR_1_2_NAND2_NUM616_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM616 (.ZN (N2014), .A1 (XNOR_1_3_NAND2_NUM616_OUT), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM617 (.ZN (N2015), .A1 (N1961), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM618_OUT, XNOR_1_2_NAND2_NUM618_OUT, XNOR_1_3_NAND2_NUM618_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM618 (.ZN (XNOR_1_1_NAND2_NUM618_OUT), .A1 (N1961), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM618 (.ZN (XNOR_1_2_NAND2_NUM618_OUT), .A1 (GND), .A2 (N1635));
      NOR2_X1 XNOR_1_3_NAND2_NUM618 (.ZN (XNOR_1_3_NAND2_NUM618_OUT), .A1 (XNOR_1_1_NAND2_NUM618_OUT), .A2 (XNOR_1_2_NAND2_NUM618_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM618 (.ZN (N2016), .A1 (XNOR_1_3_NAND2_NUM618_OUT), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM619 (.ZN (N2018), .A1 (N1965), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM620 (.ZN (N2019), .A1 (N1968), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM621_OUT, XNOR_1_2_NAND2_NUM621_OUT, XNOR_1_3_NAND2_NUM621_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM621 (.ZN (XNOR_1_1_NAND2_NUM621_OUT), .A1 (N1898), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM621 (.ZN (XNOR_1_2_NAND2_NUM621_OUT), .A1 (GND), .A2 (N1999));
      NOR2_X1 XNOR_1_3_NAND2_NUM621 (.ZN (XNOR_1_3_NAND2_NUM621_OUT), .A1 (XNOR_1_1_NAND2_NUM621_OUT), .A2 (XNOR_1_2_NAND2_NUM621_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM621 (.ZN (N2020), .A1 (XNOR_1_3_NAND2_NUM621_OUT), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM622 (.ZN (N2021), .A1 (N1987), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM623_OUT, XNOR_1_2_NAND2_NUM623_OUT, XNOR_1_3_NAND2_NUM623_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM623 (.ZN (XNOR_1_1_NAND2_NUM623_OUT), .A1 (N1987), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM623 (.ZN (XNOR_1_2_NAND2_NUM623_OUT), .A1 (GND), .A2 (N1591));
      NOR2_X1 XNOR_1_3_NAND2_NUM623 (.ZN (XNOR_1_3_NAND2_NUM623_OUT), .A1 (XNOR_1_1_NAND2_NUM623_OUT), .A2 (XNOR_1_2_NAND2_NUM623_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM623 (.ZN (N2022), .A1 (XNOR_1_3_NAND2_NUM623_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM624_OUT, XNOR_1_2_NAND2_NUM624_OUT, XNOR_1_3_NAND2_NUM624_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM624 (.ZN (XNOR_1_1_NAND2_NUM624_OUT), .A1 (N1440), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM624 (.ZN (XNOR_1_2_NAND2_NUM624_OUT), .A1 (GND), .A2 (N2002));
      NOR2_X1 XNOR_1_3_NAND2_NUM624 (.ZN (XNOR_1_3_NAND2_NUM624_OUT), .A1 (XNOR_1_1_NAND2_NUM624_OUT), .A2 (XNOR_1_2_NAND2_NUM624_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM624 (.ZN (N2023), .A1 (XNOR_1_3_NAND2_NUM624_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM625_OUT, XNOR_1_2_NAND2_NUM625_OUT, XNOR_1_3_NAND2_NUM625_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM625 (.ZN (XNOR_1_1_NAND2_NUM625_OUT), .A1 (N1261), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM625 (.ZN (XNOR_1_2_NAND2_NUM625_OUT), .A1 (GND), .A2 (N2005));
      NOR2_X1 XNOR_1_3_NAND2_NUM625 (.ZN (XNOR_1_3_NAND2_NUM625_OUT), .A1 (XNOR_1_1_NAND2_NUM625_OUT), .A2 (XNOR_1_2_NAND2_NUM625_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM625 (.ZN (N2024), .A1 (XNOR_1_3_NAND2_NUM625_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM626_OUT, XNOR_1_2_NAND2_NUM626_OUT, XNOR_1_3_NAND2_NUM626_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM626 (.ZN (XNOR_1_1_NAND2_NUM626_OUT), .A1 (N1258), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM626 (.ZN (XNOR_1_2_NAND2_NUM626_OUT), .A1 (GND), .A2 (N2007));
      NOR2_X1 XNOR_1_3_NAND2_NUM626 (.ZN (XNOR_1_3_NAND2_NUM626_OUT), .A1 (XNOR_1_1_NAND2_NUM626_OUT), .A2 (XNOR_1_2_NAND2_NUM626_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM626 (.ZN (N2025), .A1 (XNOR_1_3_NAND2_NUM626_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM627_OUT, XNOR_1_2_NAND2_NUM627_OUT, XNOR_1_3_NAND2_NUM627_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM627 (.ZN (XNOR_1_1_NAND2_NUM627_OUT), .A1 (N1975), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM627 (.ZN (XNOR_1_2_NAND2_NUM627_OUT), .A1 (GND), .A2 (N2008));
      NOR2_X1 XNOR_1_3_NAND2_NUM627 (.ZN (XNOR_1_3_NAND2_NUM627_OUT), .A1 (XNOR_1_1_NAND2_NUM627_OUT), .A2 (XNOR_1_2_NAND2_NUM627_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM627 (.ZN (N2026), .A1 (XNOR_1_3_NAND2_NUM627_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM628_OUT, XNOR_1_2_NAND2_NUM628_OUT, XNOR_1_3_NAND2_NUM628_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM628 (.ZN (XNOR_1_1_NAND2_NUM628_OUT), .A1 (N1977), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM628 (.ZN (XNOR_1_2_NAND2_NUM628_OUT), .A1 (GND), .A2 (N2009));
      NOR2_X1 XNOR_1_3_NAND2_NUM628 (.ZN (XNOR_1_3_NAND2_NUM628_OUT), .A1 (XNOR_1_1_NAND2_NUM628_OUT), .A2 (XNOR_1_2_NAND2_NUM628_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM628 (.ZN (N2027), .A1 (XNOR_1_3_NAND2_NUM628_OUT), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM629 (.ZN (N2030), .A1 (N1980), .A2 (GND));
      wire XNOR_1_1_BUFF1_NUM630_OUT;
      NOR2_X1 XNOR_1_1_BUFF1_NUM630 (.ZN (XNOR_1_1_BUFF1_NUM630_OUT), .A1 (N1980), .A2 (GND));
      NOR2_X1 XNOR_1_2_BUFF1_NUM630 (.ZN (N2033), .A1 (XNOR_1_1_BUFF1_NUM630_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM631_OUT, XNOR_1_2_NAND2_NUM631_OUT, XNOR_1_3_NAND2_NUM631_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM631 (.ZN (XNOR_1_1_NAND2_NUM631_OUT), .A1 (N1875), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM631 (.ZN (XNOR_1_2_NAND2_NUM631_OUT), .A1 (GND), .A2 (N2013));
      NOR2_X1 XNOR_1_3_NAND2_NUM631 (.ZN (XNOR_1_3_NAND2_NUM631_OUT), .A1 (XNOR_1_1_NAND2_NUM631_OUT), .A2 (XNOR_1_2_NAND2_NUM631_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM631 (.ZN (N2036), .A1 (XNOR_1_3_NAND2_NUM631_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM632_OUT, XNOR_1_2_NAND2_NUM632_OUT, XNOR_1_3_NAND2_NUM632_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM632 (.ZN (XNOR_1_1_NAND2_NUM632_OUT), .A1 (N1571), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM632 (.ZN (XNOR_1_2_NAND2_NUM632_OUT), .A1 (GND), .A2 (N2015));
      NOR2_X1 XNOR_1_3_NAND2_NUM632 (.ZN (XNOR_1_3_NAND2_NUM632_OUT), .A1 (XNOR_1_1_NAND2_NUM632_OUT), .A2 (XNOR_1_2_NAND2_NUM632_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM632 (.ZN (N2037), .A1 (XNOR_1_3_NAND2_NUM632_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM633_OUT, XNOR_1_2_NAND2_NUM633_OUT, XNOR_1_3_NAND2_NUM633_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM633 (.ZN (XNOR_1_1_NAND2_NUM633_OUT), .A1 (N2020), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM633 (.ZN (XNOR_1_2_NAND2_NUM633_OUT), .A1 (GND), .A2 (N2000));
      NOR2_X1 XNOR_1_3_NAND2_NUM633 (.ZN (XNOR_1_3_NAND2_NUM633_OUT), .A1 (XNOR_1_1_NAND2_NUM633_OUT), .A2 (XNOR_1_2_NAND2_NUM633_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM633 (.ZN (N2038), .A1 (XNOR_1_3_NAND2_NUM633_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM634_OUT, XNOR_1_2_NAND2_NUM634_OUT, XNOR_1_3_NAND2_NUM634_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM634 (.ZN (XNOR_1_1_NAND2_NUM634_OUT), .A1 (N1534), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM634 (.ZN (XNOR_1_2_NAND2_NUM634_OUT), .A1 (GND), .A2 (N2021));
      NOR2_X1 XNOR_1_3_NAND2_NUM634 (.ZN (XNOR_1_3_NAND2_NUM634_OUT), .A1 (XNOR_1_1_NAND2_NUM634_OUT), .A2 (XNOR_1_2_NAND2_NUM634_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM634 (.ZN (N2039), .A1 (XNOR_1_3_NAND2_NUM634_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM635_OUT, XNOR_1_2_NAND2_NUM635_OUT, XNOR_1_3_NAND2_NUM635_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM635 (.ZN (XNOR_1_1_NAND2_NUM635_OUT), .A1 (N2023), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM635 (.ZN (XNOR_1_2_NAND2_NUM635_OUT), .A1 (GND), .A2 (N2003));
      NOR2_X1 XNOR_1_3_NAND2_NUM635 (.ZN (XNOR_1_3_NAND2_NUM635_OUT), .A1 (XNOR_1_1_NAND2_NUM635_OUT), .A2 (XNOR_1_2_NAND2_NUM635_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM635 (.ZN (N2040), .A1 (XNOR_1_3_NAND2_NUM635_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM636_OUT, XNOR_1_2_NAND2_NUM636_OUT, XNOR_1_3_NAND2_NUM636_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM636 (.ZN (XNOR_1_1_NAND2_NUM636_OUT), .A1 (N2004), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM636 (.ZN (XNOR_1_2_NAND2_NUM636_OUT), .A1 (GND), .A2 (N2024));
      NOR2_X1 XNOR_1_3_NAND2_NUM636 (.ZN (XNOR_1_3_NAND2_NUM636_OUT), .A1 (XNOR_1_1_NAND2_NUM636_OUT), .A2 (XNOR_1_2_NAND2_NUM636_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM636 (.ZN (N2041), .A1 (XNOR_1_3_NAND2_NUM636_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM637_OUT, XNOR_1_2_NAND2_NUM637_OUT, XNOR_1_3_NAND2_NUM637_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM637 (.ZN (XNOR_1_1_NAND2_NUM637_OUT), .A1 (N2006), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM637 (.ZN (XNOR_1_2_NAND2_NUM637_OUT), .A1 (GND), .A2 (N2025));
      NOR2_X1 XNOR_1_3_NAND2_NUM637 (.ZN (XNOR_1_3_NAND2_NUM637_OUT), .A1 (XNOR_1_1_NAND2_NUM637_OUT), .A2 (XNOR_1_2_NAND2_NUM637_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM637 (.ZN (N2042), .A1 (XNOR_1_3_NAND2_NUM637_OUT), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM638 (.ZN (N2047), .A1 (N2026), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM639_OUT, XNOR_1_2_NAND2_NUM639_OUT, XNOR_1_3_NAND2_NUM639_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM639 (.ZN (XNOR_1_1_NAND2_NUM639_OUT), .A1 (N2036), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM639 (.ZN (XNOR_1_2_NAND2_NUM639_OUT), .A1 (GND), .A2 (N2014));
      NOR2_X1 XNOR_1_3_NAND2_NUM639 (.ZN (XNOR_1_3_NAND2_NUM639_OUT), .A1 (XNOR_1_1_NAND2_NUM639_OUT), .A2 (XNOR_1_2_NAND2_NUM639_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM639 (.ZN (N2052), .A1 (XNOR_1_3_NAND2_NUM639_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM640_OUT, XNOR_1_2_NAND2_NUM640_OUT, XNOR_1_3_NAND2_NUM640_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM640 (.ZN (XNOR_1_1_NAND2_NUM640_OUT), .A1 (N2037), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM640 (.ZN (XNOR_1_2_NAND2_NUM640_OUT), .A1 (GND), .A2 (N2016));
      NOR2_X1 XNOR_1_3_NAND2_NUM640 (.ZN (XNOR_1_3_NAND2_NUM640_OUT), .A1 (XNOR_1_1_NAND2_NUM640_OUT), .A2 (XNOR_1_2_NAND2_NUM640_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM640 (.ZN (N2055), .A1 (XNOR_1_3_NAND2_NUM640_OUT), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM641 (.ZN (N2060), .A1 (N2038), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM642_OUT, XNOR_1_2_NAND2_NUM642_OUT, XNOR_1_3_NAND2_NUM642_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM642 (.ZN (XNOR_1_1_NAND2_NUM642_OUT), .A1 (N2039), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM642 (.ZN (XNOR_1_2_NAND2_NUM642_OUT), .A1 (GND), .A2 (N2022));
      NOR2_X1 XNOR_1_3_NAND2_NUM642 (.ZN (XNOR_1_3_NAND2_NUM642_OUT), .A1 (XNOR_1_1_NAND2_NUM642_OUT), .A2 (XNOR_1_2_NAND2_NUM642_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM642 (.ZN (N2061), .A1 (XNOR_1_3_NAND2_NUM642_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM643_OUT, XNOR_1_2_NAND2_NUM643_OUT, XNOR_1_3_NAND2_NUM643_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM643 (.ZN (XNOR_1_1_NAND2_NUM643_OUT), .A1 (N2040), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM643 (.ZN (XNOR_1_2_NAND2_NUM643_OUT), .A1 (GND), .A2 (N290));
      NOR2_X1 XNOR_1_3_NAND2_NUM643 (.ZN (XNOR_1_3_NAND2_NUM643_OUT), .A1 (XNOR_1_1_NAND2_NUM643_OUT), .A2 (XNOR_1_2_NAND2_NUM643_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM643 (.ZN (N2062), .A1 (XNOR_1_3_NAND2_NUM643_OUT), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM644 (.ZN (N2067), .A1 (N2041), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM645 (.ZN (N2068), .A1 (N2027), .A2 (GND));
      wire XNOR_1_1_BUFF1_NUM646_OUT;
      NOR2_X1 XNOR_1_1_BUFF1_NUM646 (.ZN (XNOR_1_1_BUFF1_NUM646_OUT), .A1 (N2027), .A2 (GND));
      NOR2_X1 XNOR_1_2_BUFF1_NUM646 (.ZN (N2071), .A1 (XNOR_1_1_BUFF1_NUM646_OUT), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM647 (.ZN (N2076), .A1 (N2052), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM648 (.ZN (N2077), .A1 (N2055), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM649_OUT, XNOR_1_2_NAND2_NUM649_OUT, XNOR_1_3_NAND2_NUM649_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM649 (.ZN (XNOR_1_1_NAND2_NUM649_OUT), .A1 (N2060), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM649 (.ZN (XNOR_1_2_NAND2_NUM649_OUT), .A1 (GND), .A2 (N290));
      NOR2_X1 XNOR_1_3_NAND2_NUM649 (.ZN (XNOR_1_3_NAND2_NUM649_OUT), .A1 (XNOR_1_1_NAND2_NUM649_OUT), .A2 (XNOR_1_2_NAND2_NUM649_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM649 (.ZN (N2078), .A1 (XNOR_1_3_NAND2_NUM649_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM650_OUT, XNOR_1_2_NAND2_NUM650_OUT, XNOR_1_3_NAND2_NUM650_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM650 (.ZN (XNOR_1_1_NAND2_NUM650_OUT), .A1 (N2061), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM650 (.ZN (XNOR_1_2_NAND2_NUM650_OUT), .A1 (GND), .A2 (N290));
      NOR2_X1 XNOR_1_3_NAND2_NUM650 (.ZN (XNOR_1_3_NAND2_NUM650_OUT), .A1 (XNOR_1_1_NAND2_NUM650_OUT), .A2 (XNOR_1_2_NAND2_NUM650_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM650 (.ZN (N2081), .A1 (XNOR_1_3_NAND2_NUM650_OUT), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM651 (.ZN (N2086), .A1 (N2042), .A2 (GND));
      wire XNOR_1_1_BUFF1_NUM652_OUT;
      NOR2_X1 XNOR_1_1_BUFF1_NUM652 (.ZN (XNOR_1_1_BUFF1_NUM652_OUT), .A1 (N2042), .A2 (GND));
      NOR2_X1 XNOR_1_2_BUFF1_NUM652 (.ZN (N2089), .A1 (XNOR_1_1_BUFF1_NUM652_OUT), .A2 (GND));
      wire XNOR_1_1_AND2_NUM653_OUT, XNOR_1_2_AND2_NUM653_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM653 (.ZN (XNOR_1_1_AND2_NUM653_OUT), .A1 (N2030), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM653 (.ZN (XNOR_1_2_AND2_NUM653_OUT), .A1 (GND), .A2 (N2068));
      NOR2_X1 XNOR_1_3_AND2_NUM653 (.ZN (N2104), .A1 (XNOR_1_1_AND2_NUM653_OUT), .A2 (XNOR_1_2_AND2_NUM653_OUT));
      wire XNOR_1_1_AND2_NUM654_OUT, XNOR_1_2_AND2_NUM654_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM654 (.ZN (XNOR_1_1_AND2_NUM654_OUT), .A1 (N2033), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM654 (.ZN (XNOR_1_2_AND2_NUM654_OUT), .A1 (GND), .A2 (N2068));
      NOR2_X1 XNOR_1_3_AND2_NUM654 (.ZN (N2119), .A1 (XNOR_1_1_AND2_NUM654_OUT), .A2 (XNOR_1_2_AND2_NUM654_OUT));
      wire XNOR_1_1_AND2_NUM655_OUT, XNOR_1_2_AND2_NUM655_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM655 (.ZN (XNOR_1_1_AND2_NUM655_OUT), .A1 (N2030), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM655 (.ZN (XNOR_1_2_AND2_NUM655_OUT), .A1 (GND), .A2 (N2071));
      NOR2_X1 XNOR_1_3_AND2_NUM655 (.ZN (N2129), .A1 (XNOR_1_1_AND2_NUM655_OUT), .A2 (XNOR_1_2_AND2_NUM655_OUT));
      wire XNOR_1_1_AND2_NUM656_OUT, XNOR_1_2_AND2_NUM656_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM656 (.ZN (XNOR_1_1_AND2_NUM656_OUT), .A1 (N2033), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM656 (.ZN (XNOR_1_2_AND2_NUM656_OUT), .A1 (GND), .A2 (N2071));
      NOR2_X1 XNOR_1_3_AND2_NUM656 (.ZN (N2143), .A1 (XNOR_1_1_AND2_NUM656_OUT), .A2 (XNOR_1_2_AND2_NUM656_OUT));
      wire XNOR_1_1_BUFF1_NUM657_OUT;
      NOR2_X1 XNOR_1_1_BUFF1_NUM657 (.ZN (XNOR_1_1_BUFF1_NUM657_OUT), .A1 (N2062), .A2 (GND));
      NOR2_X1 XNOR_1_2_BUFF1_NUM657 (.ZN (N2148), .A1 (XNOR_1_1_BUFF1_NUM657_OUT), .A2 (GND));
      wire XNOR_1_1_BUFF1_NUM658_OUT;
      NOR2_X1 XNOR_1_1_BUFF1_NUM658 (.ZN (XNOR_1_1_BUFF1_NUM658_OUT), .A1 (N2062), .A2 (GND));
      NOR2_X1 XNOR_1_2_BUFF1_NUM658 (.ZN (N2151), .A1 (XNOR_1_1_BUFF1_NUM658_OUT), .A2 (GND));
      wire XNOR_1_1_BUFF1_NUM659_OUT;
      NOR2_X1 XNOR_1_1_BUFF1_NUM659 (.ZN (XNOR_1_1_BUFF1_NUM659_OUT), .A1 (N2078), .A2 (GND));
      NOR2_X1 XNOR_1_2_BUFF1_NUM659 (.ZN (N2196), .A1 (XNOR_1_1_BUFF1_NUM659_OUT), .A2 (GND));
      wire XNOR_1_1_BUFF1_NUM660_OUT;
      NOR2_X1 XNOR_1_1_BUFF1_NUM660 (.ZN (XNOR_1_1_BUFF1_NUM660_OUT), .A1 (N2078), .A2 (GND));
      NOR2_X1 XNOR_1_2_BUFF1_NUM660 (.ZN (N2199), .A1 (XNOR_1_1_BUFF1_NUM660_OUT), .A2 (GND));
      wire XNOR_1_1_BUFF1_NUM661_OUT;
      NOR2_X1 XNOR_1_1_BUFF1_NUM661 (.ZN (XNOR_1_1_BUFF1_NUM661_OUT), .A1 (N2081), .A2 (GND));
      NOR2_X1 XNOR_1_2_BUFF1_NUM661 (.ZN (N2202), .A1 (XNOR_1_1_BUFF1_NUM661_OUT), .A2 (GND));
      wire XNOR_1_1_BUFF1_NUM662_OUT;
      NOR2_X1 XNOR_1_1_BUFF1_NUM662 (.ZN (XNOR_1_1_BUFF1_NUM662_OUT), .A1 (N2081), .A2 (GND));
      NOR2_X1 XNOR_1_2_BUFF1_NUM662 (.ZN (N2205), .A1 (XNOR_1_1_BUFF1_NUM662_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM663_OUT, XNOR_1_2_NAND2_NUM663_OUT, XNOR_1_3_NAND2_NUM663_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM663 (.ZN (XNOR_1_1_NAND2_NUM663_OUT), .A1 (N2151), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM663 (.ZN (XNOR_1_2_NAND2_NUM663_OUT), .A1 (GND), .A2 (N915));
      NOR2_X1 XNOR_1_3_NAND2_NUM663 (.ZN (XNOR_1_3_NAND2_NUM663_OUT), .A1 (XNOR_1_1_NAND2_NUM663_OUT), .A2 (XNOR_1_2_NAND2_NUM663_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM663 (.ZN (N2214), .A1 (XNOR_1_3_NAND2_NUM663_OUT), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM664 (.ZN (N2215), .A1 (N2151), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM665_OUT, XNOR_1_2_NAND2_NUM665_OUT, XNOR_1_3_NAND2_NUM665_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM665 (.ZN (XNOR_1_1_NAND2_NUM665_OUT), .A1 (N2148), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM665 (.ZN (XNOR_1_2_NAND2_NUM665_OUT), .A1 (GND), .A2 (N916));
      NOR2_X1 XNOR_1_3_NAND2_NUM665 (.ZN (XNOR_1_3_NAND2_NUM665_OUT), .A1 (XNOR_1_1_NAND2_NUM665_OUT), .A2 (XNOR_1_2_NAND2_NUM665_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM665 (.ZN (N2216), .A1 (XNOR_1_3_NAND2_NUM665_OUT), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM666 (.ZN (N2217), .A1 (N2148), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM667_OUT, XNOR_1_2_NAND2_NUM667_OUT, XNOR_1_3_NAND2_NUM667_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM667 (.ZN (XNOR_1_1_NAND2_NUM667_OUT), .A1 (N2199), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM667 (.ZN (XNOR_1_2_NAND2_NUM667_OUT), .A1 (GND), .A2 (N1348));
      NOR2_X1 XNOR_1_3_NAND2_NUM667 (.ZN (XNOR_1_3_NAND2_NUM667_OUT), .A1 (XNOR_1_1_NAND2_NUM667_OUT), .A2 (XNOR_1_2_NAND2_NUM667_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM667 (.ZN (N2222), .A1 (XNOR_1_3_NAND2_NUM667_OUT), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM668 (.ZN (N2223), .A1 (N2199), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM669_OUT, XNOR_1_2_NAND2_NUM669_OUT, XNOR_1_3_NAND2_NUM669_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM669 (.ZN (XNOR_1_1_NAND2_NUM669_OUT), .A1 (N2196), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM669 (.ZN (XNOR_1_2_NAND2_NUM669_OUT), .A1 (GND), .A2 (N1349));
      NOR2_X1 XNOR_1_3_NAND2_NUM669 (.ZN (XNOR_1_3_NAND2_NUM669_OUT), .A1 (XNOR_1_1_NAND2_NUM669_OUT), .A2 (XNOR_1_2_NAND2_NUM669_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM669 (.ZN (N2224), .A1 (XNOR_1_3_NAND2_NUM669_OUT), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM670 (.ZN (N2225), .A1 (N2196), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM671_OUT, XNOR_1_2_NAND2_NUM671_OUT, XNOR_1_3_NAND2_NUM671_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM671 (.ZN (XNOR_1_1_NAND2_NUM671_OUT), .A1 (N2205), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM671 (.ZN (XNOR_1_2_NAND2_NUM671_OUT), .A1 (GND), .A2 (N913));
      NOR2_X1 XNOR_1_3_NAND2_NUM671 (.ZN (XNOR_1_3_NAND2_NUM671_OUT), .A1 (XNOR_1_1_NAND2_NUM671_OUT), .A2 (XNOR_1_2_NAND2_NUM671_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM671 (.ZN (N2226), .A1 (XNOR_1_3_NAND2_NUM671_OUT), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM672 (.ZN (N2227), .A1 (N2205), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM673_OUT, XNOR_1_2_NAND2_NUM673_OUT, XNOR_1_3_NAND2_NUM673_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM673 (.ZN (XNOR_1_1_NAND2_NUM673_OUT), .A1 (N2202), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM673 (.ZN (XNOR_1_2_NAND2_NUM673_OUT), .A1 (GND), .A2 (N914));
      NOR2_X1 XNOR_1_3_NAND2_NUM673 (.ZN (XNOR_1_3_NAND2_NUM673_OUT), .A1 (XNOR_1_1_NAND2_NUM673_OUT), .A2 (XNOR_1_2_NAND2_NUM673_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM673 (.ZN (N2228), .A1 (XNOR_1_3_NAND2_NUM673_OUT), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM674 (.ZN (N2229), .A1 (N2202), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM675_OUT, XNOR_1_2_NAND2_NUM675_OUT, XNOR_1_3_NAND2_NUM675_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM675 (.ZN (XNOR_1_1_NAND2_NUM675_OUT), .A1 (N667), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM675 (.ZN (XNOR_1_2_NAND2_NUM675_OUT), .A1 (GND), .A2 (N2215));
      NOR2_X1 XNOR_1_3_NAND2_NUM675 (.ZN (XNOR_1_3_NAND2_NUM675_OUT), .A1 (XNOR_1_1_NAND2_NUM675_OUT), .A2 (XNOR_1_2_NAND2_NUM675_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM675 (.ZN (N2230), .A1 (XNOR_1_3_NAND2_NUM675_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM676_OUT, XNOR_1_2_NAND2_NUM676_OUT, XNOR_1_3_NAND2_NUM676_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM676 (.ZN (XNOR_1_1_NAND2_NUM676_OUT), .A1 (N664), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM676 (.ZN (XNOR_1_2_NAND2_NUM676_OUT), .A1 (GND), .A2 (N2217));
      NOR2_X1 XNOR_1_3_NAND2_NUM676 (.ZN (XNOR_1_3_NAND2_NUM676_OUT), .A1 (XNOR_1_1_NAND2_NUM676_OUT), .A2 (XNOR_1_2_NAND2_NUM676_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM676 (.ZN (N2231), .A1 (XNOR_1_3_NAND2_NUM676_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM677_OUT, XNOR_1_2_NAND2_NUM677_OUT, XNOR_1_3_NAND2_NUM677_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM677 (.ZN (XNOR_1_1_NAND2_NUM677_OUT), .A1 (N1255), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM677 (.ZN (XNOR_1_2_NAND2_NUM677_OUT), .A1 (GND), .A2 (N2223));
      NOR2_X1 XNOR_1_3_NAND2_NUM677 (.ZN (XNOR_1_3_NAND2_NUM677_OUT), .A1 (XNOR_1_1_NAND2_NUM677_OUT), .A2 (XNOR_1_2_NAND2_NUM677_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM677 (.ZN (N2232), .A1 (XNOR_1_3_NAND2_NUM677_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM678_OUT, XNOR_1_2_NAND2_NUM678_OUT, XNOR_1_3_NAND2_NUM678_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM678 (.ZN (XNOR_1_1_NAND2_NUM678_OUT), .A1 (N1252), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM678 (.ZN (XNOR_1_2_NAND2_NUM678_OUT), .A1 (GND), .A2 (N2225));
      NOR2_X1 XNOR_1_3_NAND2_NUM678 (.ZN (XNOR_1_3_NAND2_NUM678_OUT), .A1 (XNOR_1_1_NAND2_NUM678_OUT), .A2 (XNOR_1_2_NAND2_NUM678_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM678 (.ZN (N2233), .A1 (XNOR_1_3_NAND2_NUM678_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM679_OUT, XNOR_1_2_NAND2_NUM679_OUT, XNOR_1_3_NAND2_NUM679_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM679 (.ZN (XNOR_1_1_NAND2_NUM679_OUT), .A1 (N661), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM679 (.ZN (XNOR_1_2_NAND2_NUM679_OUT), .A1 (GND), .A2 (N2227));
      NOR2_X1 XNOR_1_3_NAND2_NUM679 (.ZN (XNOR_1_3_NAND2_NUM679_OUT), .A1 (XNOR_1_1_NAND2_NUM679_OUT), .A2 (XNOR_1_2_NAND2_NUM679_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM679 (.ZN (N2234), .A1 (XNOR_1_3_NAND2_NUM679_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM680_OUT, XNOR_1_2_NAND2_NUM680_OUT, XNOR_1_3_NAND2_NUM680_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM680 (.ZN (XNOR_1_1_NAND2_NUM680_OUT), .A1 (N658), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM680 (.ZN (XNOR_1_2_NAND2_NUM680_OUT), .A1 (GND), .A2 (N2229));
      NOR2_X1 XNOR_1_3_NAND2_NUM680 (.ZN (XNOR_1_3_NAND2_NUM680_OUT), .A1 (XNOR_1_1_NAND2_NUM680_OUT), .A2 (XNOR_1_2_NAND2_NUM680_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM680 (.ZN (N2235), .A1 (XNOR_1_3_NAND2_NUM680_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM681_OUT, XNOR_1_2_NAND2_NUM681_OUT, XNOR_1_3_NAND2_NUM681_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM681 (.ZN (XNOR_1_1_NAND2_NUM681_OUT), .A1 (N2214), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM681 (.ZN (XNOR_1_2_NAND2_NUM681_OUT), .A1 (GND), .A2 (N2230));
      NOR2_X1 XNOR_1_3_NAND2_NUM681 (.ZN (XNOR_1_3_NAND2_NUM681_OUT), .A1 (XNOR_1_1_NAND2_NUM681_OUT), .A2 (XNOR_1_2_NAND2_NUM681_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM681 (.ZN (N2236), .A1 (XNOR_1_3_NAND2_NUM681_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM682_OUT, XNOR_1_2_NAND2_NUM682_OUT, XNOR_1_3_NAND2_NUM682_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM682 (.ZN (XNOR_1_1_NAND2_NUM682_OUT), .A1 (N2216), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM682 (.ZN (XNOR_1_2_NAND2_NUM682_OUT), .A1 (GND), .A2 (N2231));
      NOR2_X1 XNOR_1_3_NAND2_NUM682 (.ZN (XNOR_1_3_NAND2_NUM682_OUT), .A1 (XNOR_1_1_NAND2_NUM682_OUT), .A2 (XNOR_1_2_NAND2_NUM682_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM682 (.ZN (N2237), .A1 (XNOR_1_3_NAND2_NUM682_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM683_OUT, XNOR_1_2_NAND2_NUM683_OUT, XNOR_1_3_NAND2_NUM683_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM683 (.ZN (XNOR_1_1_NAND2_NUM683_OUT), .A1 (N2222), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM683 (.ZN (XNOR_1_2_NAND2_NUM683_OUT), .A1 (GND), .A2 (N2232));
      NOR2_X1 XNOR_1_3_NAND2_NUM683 (.ZN (XNOR_1_3_NAND2_NUM683_OUT), .A1 (XNOR_1_1_NAND2_NUM683_OUT), .A2 (XNOR_1_2_NAND2_NUM683_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM683 (.ZN (N2240), .A1 (XNOR_1_3_NAND2_NUM683_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM684_OUT, XNOR_1_2_NAND2_NUM684_OUT, XNOR_1_3_NAND2_NUM684_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM684 (.ZN (XNOR_1_1_NAND2_NUM684_OUT), .A1 (N2224), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM684 (.ZN (XNOR_1_2_NAND2_NUM684_OUT), .A1 (GND), .A2 (N2233));
      NOR2_X1 XNOR_1_3_NAND2_NUM684 (.ZN (XNOR_1_3_NAND2_NUM684_OUT), .A1 (XNOR_1_1_NAND2_NUM684_OUT), .A2 (XNOR_1_2_NAND2_NUM684_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM684 (.ZN (N2241), .A1 (XNOR_1_3_NAND2_NUM684_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM685_OUT, XNOR_1_2_NAND2_NUM685_OUT, XNOR_1_3_NAND2_NUM685_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM685 (.ZN (XNOR_1_1_NAND2_NUM685_OUT), .A1 (N2226), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM685 (.ZN (XNOR_1_2_NAND2_NUM685_OUT), .A1 (GND), .A2 (N2234));
      NOR2_X1 XNOR_1_3_NAND2_NUM685 (.ZN (XNOR_1_3_NAND2_NUM685_OUT), .A1 (XNOR_1_1_NAND2_NUM685_OUT), .A2 (XNOR_1_2_NAND2_NUM685_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM685 (.ZN (N2244), .A1 (XNOR_1_3_NAND2_NUM685_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM686_OUT, XNOR_1_2_NAND2_NUM686_OUT, XNOR_1_3_NAND2_NUM686_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM686 (.ZN (XNOR_1_1_NAND2_NUM686_OUT), .A1 (N2228), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM686 (.ZN (XNOR_1_2_NAND2_NUM686_OUT), .A1 (GND), .A2 (N2235));
      NOR2_X1 XNOR_1_3_NAND2_NUM686 (.ZN (XNOR_1_3_NAND2_NUM686_OUT), .A1 (XNOR_1_1_NAND2_NUM686_OUT), .A2 (XNOR_1_2_NAND2_NUM686_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM686 (.ZN (N2245), .A1 (XNOR_1_3_NAND2_NUM686_OUT), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM687 (.ZN (N2250), .A1 (N2236), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM688 (.ZN (N2253), .A1 (N2240), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM689 (.ZN (N2256), .A1 (N2244), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM690 (.ZN (N2257), .A1 (N2237), .A2 (GND));
      wire XNOR_1_1_BUFF1_NUM691_OUT;
      NOR2_X1 XNOR_1_1_BUFF1_NUM691 (.ZN (XNOR_1_1_BUFF1_NUM691_OUT), .A1 (N2237), .A2 (GND));
      NOR2_X1 XNOR_1_2_BUFF1_NUM691 (.ZN (N2260), .A1 (XNOR_1_1_BUFF1_NUM691_OUT), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM692 (.ZN (N2263), .A1 (N2241), .A2 (GND));
      wire XNOR_1_1_AND2_NUM693_OUT, XNOR_1_2_AND2_NUM693_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM693 (.ZN (XNOR_1_1_AND2_NUM693_OUT), .A1 (N1164), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM693 (.ZN (XNOR_1_2_AND2_NUM693_OUT), .A1 (GND), .A2 (N2241));
      NOR2_X1 XNOR_1_3_AND2_NUM693 (.ZN (N2266), .A1 (XNOR_1_1_AND2_NUM693_OUT), .A2 (XNOR_1_2_AND2_NUM693_OUT));
      NOR2_X1 XNOR_NOT1_NUM694 (.ZN (N2269), .A1 (N2245), .A2 (GND));
      wire XNOR_1_1_AND2_NUM695_OUT, XNOR_1_2_AND2_NUM695_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM695 (.ZN (XNOR_1_1_AND2_NUM695_OUT), .A1 (N1168), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM695 (.ZN (XNOR_1_2_AND2_NUM695_OUT), .A1 (GND), .A2 (N2245));
      NOR2_X1 XNOR_1_3_AND2_NUM695 (.ZN (N2272), .A1 (XNOR_1_1_AND2_NUM695_OUT), .A2 (XNOR_1_2_AND2_NUM695_OUT));
      wire XNOR_1_1_NAND8_NUM696_OUT, XNOR_1_2_NAND8_NUM696_OUT, XNOR_1_3_NAND8_NUM696_OUT;
      NOR2_X1 XNOR_1_1_NAND8_NUM696 (.ZN (XNOR_1_1_NAND8_NUM696_OUT), .A1 (N2067), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND8_NUM696 (.ZN (XNOR_1_2_NAND8_NUM696_OUT), .A1 (GND), .A2 (N2012));
      NOR2_X1 XNOR_1_3_NAND8_NUM696 (.ZN (XNOR_1_3_NAND8_NUM696_OUT), .A1 (XNOR_1_1_NAND8_NUM696_OUT), .A2 (XNOR_1_2_NAND8_NUM696_OUT));

      wire XNOR_2_1_NAND8_NUM696_OUT, XNOR_2_2_NAND8_NUM696_OUT, XNOR_2_3_NAND8_NUM696_OUT;
      NOR2_X1 XNOR_2_1_NAND8_NUM696 (.ZN (XNOR_2_1_NAND8_NUM696_OUT), .A1 (N2047), .A2 (GND));
      NOR2_X1 XNOR_2_2_NAND8_NUM696 (.ZN (XNOR_2_2_NAND8_NUM696_OUT), .A1 (GND), .A2 (N2250));
      NOR2_X1 XNOR_2_3_NAND8_NUM696 (.ZN (XNOR_2_3_NAND8_NUM696_OUT), .A1 (XNOR_2_1_NAND8_NUM696_OUT), .A2 (XNOR_2_2_NAND8_NUM696_OUT));

      wire XNOR_3_1_NAND8_NUM696_OUT, XNOR_3_2_NAND8_NUM696_OUT, XNOR_3_3_NAND8_NUM696_OUT;
      NOR2_X1 XNOR_3_1_NAND8_NUM696 (.ZN (XNOR_3_1_NAND8_NUM696_OUT), .A1 (N899), .A2 (GND));
      NOR2_X1 XNOR_3_2_NAND8_NUM696 (.ZN (XNOR_3_2_NAND8_NUM696_OUT), .A1 (GND), .A2 (N2256));
      NOR2_X1 XNOR_3_3_NAND8_NUM696 (.ZN (XNOR_3_3_NAND8_NUM696_OUT), .A1 (XNOR_3_1_NAND8_NUM696_OUT), .A2 (XNOR_3_2_NAND8_NUM696_OUT));

      wire XNOR_4_1_NAND8_NUM696_OUT, XNOR_4_2_NAND8_NUM696_OUT, XNOR_4_3_NAND8_NUM696_OUT;
      NOR2_X1 XNOR_4_1_NAND8_NUM696 (.ZN (XNOR_4_1_NAND8_NUM696_OUT), .A1 (N2253), .A2 (GND));
      NOR2_X1 XNOR_4_2_NAND8_NUM696 (.ZN (XNOR_4_2_NAND8_NUM696_OUT), .A1 (GND), .A2 (N903));
      NOR2_X1 XNOR_4_3_NAND8_NUM696 (.ZN (XNOR_4_3_NAND8_NUM696_OUT), .A1 (XNOR_4_1_NAND8_NUM696_OUT), .A2 (XNOR_4_2_NAND8_NUM696_OUT));

      wire XNOR_5_1_NAND8_NUM696_OUT, XNOR_5_2_NAND8_NUM696_OUT, XNOR_5_3_NAND8_NUM696_OUT;
      NOR2_X1 XNOR_5_1_NAND8_NUM696 (.ZN (XNOR_5_1_NAND8_NUM696_OUT), .A1 (XNOR_1_3_NAND8_NUM696_OUT), .A2 (GND));
      NOR2_X1 XNOR_5_2_NAND8_NUM696 (.ZN (XNOR_5_2_NAND8_NUM696_OUT), .A1 (GND), .A2 (XNOR_2_3_NAND8_NUM696_OUT));
      NOR2_X1 XNOR_5_3_NAND8_NUM696 (.ZN (XNOR_5_3_NAND8_NUM696_OUT), .A1 (XNOR_5_1_NAND8_NUM696_OUT), .A2 (XNOR_5_2_NAND8_NUM696_OUT));

      wire XNOR_6_1_NAND8_NUM696_OUT, XNOR_6_2_NAND8_NUM696_OUT, XNOR_6_3_NAND8_NUM696_OUT;
      NOR2_X1 XNOR_6_1_NAND8_NUM696 (.ZN (XNOR_6_1_NAND8_NUM696_OUT), .A1 (XNOR_3_3_NAND8_NUM696_OUT), .A2 (GND));
      NOR2_X1 XNOR_6_2_NAND8_NUM696 (.ZN (XNOR_6_2_NAND8_NUM696_OUT), .A1 (GND), .A2 (XNOR_4_3_NAND8_NUM696_OUT));
      NOR2_X1 XNOR_6_3_NAND8_NUM696 (.ZN (XNOR_6_3_NAND8_NUM696_OUT), .A1 (XNOR_6_1_NAND8_NUM696_OUT), .A2 (XNOR_6_2_NAND8_NUM696_OUT));

      wire XNOR_7_1_NAND8_NUM696_OUT, XNOR_7_2_NAND8_NUM696_OUT, XNOR_7_3_NAND8_NUM696_OUT;
      NOR2_X1 XNOR_7_1_NAND8_NUM696 (.ZN (XNOR_7_1_NAND8_NUM696_OUT), .A1 (XNOR_5_3_NAND8_NUM696_OUT), .A2 (GND));
      NOR2_X1 XNOR_7_2_NAND8_NUM696 (.ZN (XNOR_7_2_NAND8_NUM696_OUT), .A1 (GND), .A2 (XNOR_6_3_NAND8_NUM696_OUT));
      NOR2_X1 XNOR_7_3_NAND8_NUM696 (.ZN (XNOR_7_3_NAND8_NUM696_OUT), .A1 (XNOR_7_1_NAND8_NUM696_OUT), .A2 (XNOR_7_2_NAND8_NUM696_OUT));

      NOR2_X1 XNOR_8_1_NAND8_NUM696 (.ZN (N2279), .A1 (XNOR_7_3_NAND8_NUM696_OUT), .A2 (GND));
      wire XNOR_1_1_BUFF1_NUM697_OUT;
      NOR2_X1 XNOR_1_1_BUFF1_NUM697 (.ZN (XNOR_1_1_BUFF1_NUM697_OUT), .A1 (N2266), .A2 (GND));
      NOR2_X1 XNOR_1_2_BUFF1_NUM697 (.ZN (N2286), .A1 (XNOR_1_1_BUFF1_NUM697_OUT), .A2 (GND));
      wire XNOR_1_1_BUFF1_NUM698_OUT;
      NOR2_X1 XNOR_1_1_BUFF1_NUM698 (.ZN (XNOR_1_1_BUFF1_NUM698_OUT), .A1 (N2266), .A2 (GND));
      NOR2_X1 XNOR_1_2_BUFF1_NUM698 (.ZN (N2297), .A1 (XNOR_1_1_BUFF1_NUM698_OUT), .A2 (GND));
      wire XNOR_1_1_BUFF1_NUM699_OUT;
      NOR2_X1 XNOR_1_1_BUFF1_NUM699 (.ZN (XNOR_1_1_BUFF1_NUM699_OUT), .A1 (N2272), .A2 (GND));
      NOR2_X1 XNOR_1_2_BUFF1_NUM699 (.ZN (N2315), .A1 (XNOR_1_1_BUFF1_NUM699_OUT), .A2 (GND));
      wire XNOR_1_1_BUFF1_NUM700_OUT;
      NOR2_X1 XNOR_1_1_BUFF1_NUM700 (.ZN (XNOR_1_1_BUFF1_NUM700_OUT), .A1 (N2272), .A2 (GND));
      NOR2_X1 XNOR_1_2_BUFF1_NUM700 (.ZN (N2326), .A1 (XNOR_1_1_BUFF1_NUM700_OUT), .A2 (GND));
      wire XNOR_1_1_AND2_NUM701_OUT, XNOR_1_2_AND2_NUM701_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM701 (.ZN (XNOR_1_1_AND2_NUM701_OUT), .A1 (N2086), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM701 (.ZN (XNOR_1_2_AND2_NUM701_OUT), .A1 (GND), .A2 (N2257));
      NOR2_X1 XNOR_1_3_AND2_NUM701 (.ZN (N2340), .A1 (XNOR_1_1_AND2_NUM701_OUT), .A2 (XNOR_1_2_AND2_NUM701_OUT));
      wire XNOR_1_1_AND2_NUM702_OUT, XNOR_1_2_AND2_NUM702_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM702 (.ZN (XNOR_1_1_AND2_NUM702_OUT), .A1 (N2089), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM702 (.ZN (XNOR_1_2_AND2_NUM702_OUT), .A1 (GND), .A2 (N2257));
      NOR2_X1 XNOR_1_3_AND2_NUM702 (.ZN (N2353), .A1 (XNOR_1_1_AND2_NUM702_OUT), .A2 (XNOR_1_2_AND2_NUM702_OUT));
      wire XNOR_1_1_AND2_NUM703_OUT, XNOR_1_2_AND2_NUM703_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM703 (.ZN (XNOR_1_1_AND2_NUM703_OUT), .A1 (N2086), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM703 (.ZN (XNOR_1_2_AND2_NUM703_OUT), .A1 (GND), .A2 (N2260));
      NOR2_X1 XNOR_1_3_AND2_NUM703 (.ZN (N2361), .A1 (XNOR_1_1_AND2_NUM703_OUT), .A2 (XNOR_1_2_AND2_NUM703_OUT));
      wire XNOR_1_1_AND2_NUM704_OUT, XNOR_1_2_AND2_NUM704_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM704 (.ZN (XNOR_1_1_AND2_NUM704_OUT), .A1 (N2089), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM704 (.ZN (XNOR_1_2_AND2_NUM704_OUT), .A1 (GND), .A2 (N2260));
      NOR2_X1 XNOR_1_3_AND2_NUM704 (.ZN (N2375), .A1 (XNOR_1_1_AND2_NUM704_OUT), .A2 (XNOR_1_2_AND2_NUM704_OUT));
      wire XNOR_1_1_AND4_NUM705_OUT, XNOR_1_2_AND4_NUM705_OUT, XNOR_1_3_AND4_NUM705_OUT;
      NOR2_X1 XNOR_1_1_AND4_NUM705 (.ZN (XNOR_1_1_AND4_NUM705_OUT), .A1 (N338), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND4_NUM705 (.ZN (XNOR_1_2_AND4_NUM705_OUT), .A1 (GND), .A2 (N2279));
      NOR2_X1 XNOR_1_3_AND4_NUM705 (.ZN (XNOR_1_3_AND4_NUM705_OUT), .A1 (XNOR_1_1_AND4_NUM705_OUT), .A2 (XNOR_1_2_AND4_NUM705_OUT));

      wire XNOR_2_1_AND4_NUM705_OUT, XNOR_2_2_AND4_NUM705_OUT, XNOR_2_3_AND4_NUM705_OUT;
      NOR2_X1 XNOR_2_1_AND4_NUM705 (.ZN (XNOR_2_1_AND4_NUM705_OUT), .A1 (N313), .A2 (GND));
      NOR2_X1 XNOR_2_2_AND4_NUM705 (.ZN (XNOR_2_2_AND4_NUM705_OUT), .A1 (GND), .A2 (N313));
      NOR2_X1 XNOR_2_3_AND4_NUM705 (.ZN (XNOR_2_3_AND4_NUM705_OUT), .A1 (XNOR_2_1_AND4_NUM705_OUT), .A2 (XNOR_2_2_AND4_NUM705_OUT));

      wire XNOR_3_1_AND4_NUM705_OUT, XNOR_3_2_AND4_NUM705_OUT;
      NOR2_X1 XNOR_3_1_AND4_NUM705 (.ZN (XNOR_3_1_AND4_NUM705_OUT), .A1 (XNOR_1_3_AND4_NUM705_OUT), .A2 (GND));
      NOR2_X1 XNOR_3_2_AND4_NUM705 (.ZN (XNOR_3_2_AND4_NUM705_OUT), .A1 (GND), .A2 (XNOR_2_3_AND4_NUM705_OUT));
      NOR2_X1 XNOR_3_3_AND4_NUM705 (.ZN (N2384), .A1 (XNOR_3_1_AND4_NUM705_OUT), .A2 (XNOR_3_2_AND4_NUM705_OUT));
      wire XNOR_1_1_AND2_NUM706_OUT, XNOR_1_2_AND2_NUM706_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM706 (.ZN (XNOR_1_1_AND2_NUM706_OUT), .A1 (N1163), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM706 (.ZN (XNOR_1_2_AND2_NUM706_OUT), .A1 (GND), .A2 (N2263));
      NOR2_X1 XNOR_1_3_AND2_NUM706 (.ZN (N2385), .A1 (XNOR_1_1_AND2_NUM706_OUT), .A2 (XNOR_1_2_AND2_NUM706_OUT));
      wire XNOR_1_1_AND2_NUM707_OUT, XNOR_1_2_AND2_NUM707_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM707 (.ZN (XNOR_1_1_AND2_NUM707_OUT), .A1 (N1164), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM707 (.ZN (XNOR_1_2_AND2_NUM707_OUT), .A1 (GND), .A2 (N2263));
      NOR2_X1 XNOR_1_3_AND2_NUM707 (.ZN (N2386), .A1 (XNOR_1_1_AND2_NUM707_OUT), .A2 (XNOR_1_2_AND2_NUM707_OUT));
      wire XNOR_1_1_AND2_NUM708_OUT, XNOR_1_2_AND2_NUM708_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM708 (.ZN (XNOR_1_1_AND2_NUM708_OUT), .A1 (N1167), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM708 (.ZN (XNOR_1_2_AND2_NUM708_OUT), .A1 (GND), .A2 (N2269));
      NOR2_X1 XNOR_1_3_AND2_NUM708 (.ZN (N2426), .A1 (XNOR_1_1_AND2_NUM708_OUT), .A2 (XNOR_1_2_AND2_NUM708_OUT));
      wire XNOR_1_1_AND2_NUM709_OUT, XNOR_1_2_AND2_NUM709_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM709 (.ZN (XNOR_1_1_AND2_NUM709_OUT), .A1 (N1168), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM709 (.ZN (XNOR_1_2_AND2_NUM709_OUT), .A1 (GND), .A2 (N2269));
      NOR2_X1 XNOR_1_3_AND2_NUM709 (.ZN (N2427), .A1 (XNOR_1_1_AND2_NUM709_OUT), .A2 (XNOR_1_2_AND2_NUM709_OUT));
      wire XNOR_1_1_NAND5_NUM710_OUT, XNOR_1_2_NAND5_NUM710_OUT, XNOR_1_3_NAND5_NUM710_OUT;
      NOR2_X1 XNOR_1_1_NAND5_NUM710 (.ZN (XNOR_1_1_NAND5_NUM710_OUT), .A1 (N2286), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND5_NUM710 (.ZN (XNOR_1_2_NAND5_NUM710_OUT), .A1 (GND), .A2 (N2315));
      NOR2_X1 XNOR_1_3_NAND5_NUM710 (.ZN (XNOR_1_3_NAND5_NUM710_OUT), .A1 (XNOR_1_1_NAND5_NUM710_OUT), .A2 (XNOR_1_2_NAND5_NUM710_OUT));

      wire XNOR_2_1_NAND5_NUM710_OUT, XNOR_2_2_NAND5_NUM710_OUT, XNOR_2_3_NAND5_NUM710_OUT;
      NOR2_X1 XNOR_2_1_NAND5_NUM710 (.ZN (XNOR_2_1_NAND5_NUM710_OUT), .A1 (N2361), .A2 (GND));
      NOR2_X1 XNOR_2_2_NAND5_NUM710 (.ZN (XNOR_2_2_NAND5_NUM710_OUT), .A1 (GND), .A2 (N2104));
      NOR2_X1 XNOR_2_3_NAND5_NUM710 (.ZN (XNOR_2_3_NAND5_NUM710_OUT), .A1 (XNOR_2_1_NAND5_NUM710_OUT), .A2 (XNOR_2_2_NAND5_NUM710_OUT));

      wire XNOR_3_1_NAND5_NUM710_OUT, XNOR_3_2_NAND5_NUM710_OUT, XNOR_3_3_NAND5_NUM710_OUT;
      NOR2_X1 XNOR_3_1_NAND5_NUM710 (.ZN (XNOR_3_1_NAND5_NUM710_OUT), .A1 (XNOR_1_3_NAND5_NUM710_OUT), .A2 (GND));
      NOR2_X1 XNOR_3_2_NAND5_NUM710 (.ZN (XNOR_3_2_NAND5_NUM710_OUT), .A1 (GND), .A2 (XNOR_2_3_NAND5_NUM710_OUT));
      NOR2_X1 XNOR_3_3_NAND5_NUM710 (.ZN (XNOR_3_3_NAND5_NUM710_OUT), .A1 (XNOR_3_1_NAND5_NUM710_OUT), .A2 (XNOR_3_2_NAND5_NUM710_OUT));

      wire XNOR_4_1_NAND5_NUM710_OUT, XNOR_4_2_NAND5_NUM710_OUT, XNOR_4_3_NAND5_NUM710_OUT;
      NOR2_X1 XNOR_4_1_NAND5_NUM710 (.ZN (XNOR_4_1_NAND5_NUM710_OUT), .A1 (N1171), .A2 (GND));
      NOR2_X1 XNOR_4_2_NAND5_NUM710 (.ZN (XNOR_4_2_NAND5_NUM710_OUT), .A1 (GND), .A2 (XNOR_3_3_NAND5_NUM710_OUT));
      NOR2_X1 XNOR_4_3_NAND5_NUM710 (.ZN (XNOR_4_3_NAND5_NUM710_OUT), .A1 (XNOR_4_1_NAND5_NUM710_OUT), .A2 (XNOR_4_2_NAND5_NUM710_OUT));

      NOR2_X1 XNOR_5_1_NAND5_NUM710 (.ZN (N2537), .A1 (XNOR_4_3_NAND5_NUM710_OUT), .A2 (GND));
      wire XNOR_1_1_NAND5_NUM711_OUT, XNOR_1_2_NAND5_NUM711_OUT, XNOR_1_3_NAND5_NUM711_OUT;
      NOR2_X1 XNOR_1_1_NAND5_NUM711 (.ZN (XNOR_1_1_NAND5_NUM711_OUT), .A1 (N2286), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND5_NUM711 (.ZN (XNOR_1_2_NAND5_NUM711_OUT), .A1 (GND), .A2 (N2315));
      NOR2_X1 XNOR_1_3_NAND5_NUM711 (.ZN (XNOR_1_3_NAND5_NUM711_OUT), .A1 (XNOR_1_1_NAND5_NUM711_OUT), .A2 (XNOR_1_2_NAND5_NUM711_OUT));

      wire XNOR_2_1_NAND5_NUM711_OUT, XNOR_2_2_NAND5_NUM711_OUT, XNOR_2_3_NAND5_NUM711_OUT;
      NOR2_X1 XNOR_2_1_NAND5_NUM711 (.ZN (XNOR_2_1_NAND5_NUM711_OUT), .A1 (N2340), .A2 (GND));
      NOR2_X1 XNOR_2_2_NAND5_NUM711 (.ZN (XNOR_2_2_NAND5_NUM711_OUT), .A1 (GND), .A2 (N2129));
      NOR2_X1 XNOR_2_3_NAND5_NUM711 (.ZN (XNOR_2_3_NAND5_NUM711_OUT), .A1 (XNOR_2_1_NAND5_NUM711_OUT), .A2 (XNOR_2_2_NAND5_NUM711_OUT));

      wire XNOR_3_1_NAND5_NUM711_OUT, XNOR_3_2_NAND5_NUM711_OUT, XNOR_3_3_NAND5_NUM711_OUT;
      NOR2_X1 XNOR_3_1_NAND5_NUM711 (.ZN (XNOR_3_1_NAND5_NUM711_OUT), .A1 (XNOR_1_3_NAND5_NUM711_OUT), .A2 (GND));
      NOR2_X1 XNOR_3_2_NAND5_NUM711 (.ZN (XNOR_3_2_NAND5_NUM711_OUT), .A1 (GND), .A2 (XNOR_2_3_NAND5_NUM711_OUT));
      NOR2_X1 XNOR_3_3_NAND5_NUM711 (.ZN (XNOR_3_3_NAND5_NUM711_OUT), .A1 (XNOR_3_1_NAND5_NUM711_OUT), .A2 (XNOR_3_2_NAND5_NUM711_OUT));

      wire XNOR_4_1_NAND5_NUM711_OUT, XNOR_4_2_NAND5_NUM711_OUT, XNOR_4_3_NAND5_NUM711_OUT;
      NOR2_X1 XNOR_4_1_NAND5_NUM711 (.ZN (XNOR_4_1_NAND5_NUM711_OUT), .A1 (N1171), .A2 (GND));
      NOR2_X1 XNOR_4_2_NAND5_NUM711 (.ZN (XNOR_4_2_NAND5_NUM711_OUT), .A1 (GND), .A2 (XNOR_3_3_NAND5_NUM711_OUT));
      NOR2_X1 XNOR_4_3_NAND5_NUM711 (.ZN (XNOR_4_3_NAND5_NUM711_OUT), .A1 (XNOR_4_1_NAND5_NUM711_OUT), .A2 (XNOR_4_2_NAND5_NUM711_OUT));

      NOR2_X1 XNOR_5_1_NAND5_NUM711 (.ZN (N2540), .A1 (XNOR_4_3_NAND5_NUM711_OUT), .A2 (GND));
      wire XNOR_1_1_NAND5_NUM712_OUT, XNOR_1_2_NAND5_NUM712_OUT, XNOR_1_3_NAND5_NUM712_OUT;
      NOR2_X1 XNOR_1_1_NAND5_NUM712 (.ZN (XNOR_1_1_NAND5_NUM712_OUT), .A1 (N2286), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND5_NUM712 (.ZN (XNOR_1_2_NAND5_NUM712_OUT), .A1 (GND), .A2 (N2315));
      NOR2_X1 XNOR_1_3_NAND5_NUM712 (.ZN (XNOR_1_3_NAND5_NUM712_OUT), .A1 (XNOR_1_1_NAND5_NUM712_OUT), .A2 (XNOR_1_2_NAND5_NUM712_OUT));

      wire XNOR_2_1_NAND5_NUM712_OUT, XNOR_2_2_NAND5_NUM712_OUT, XNOR_2_3_NAND5_NUM712_OUT;
      NOR2_X1 XNOR_2_1_NAND5_NUM712 (.ZN (XNOR_2_1_NAND5_NUM712_OUT), .A1 (N2340), .A2 (GND));
      NOR2_X1 XNOR_2_2_NAND5_NUM712 (.ZN (XNOR_2_2_NAND5_NUM712_OUT), .A1 (GND), .A2 (N2119));
      NOR2_X1 XNOR_2_3_NAND5_NUM712 (.ZN (XNOR_2_3_NAND5_NUM712_OUT), .A1 (XNOR_2_1_NAND5_NUM712_OUT), .A2 (XNOR_2_2_NAND5_NUM712_OUT));

      wire XNOR_3_1_NAND5_NUM712_OUT, XNOR_3_2_NAND5_NUM712_OUT, XNOR_3_3_NAND5_NUM712_OUT;
      NOR2_X1 XNOR_3_1_NAND5_NUM712 (.ZN (XNOR_3_1_NAND5_NUM712_OUT), .A1 (XNOR_1_3_NAND5_NUM712_OUT), .A2 (GND));
      NOR2_X1 XNOR_3_2_NAND5_NUM712 (.ZN (XNOR_3_2_NAND5_NUM712_OUT), .A1 (GND), .A2 (XNOR_2_3_NAND5_NUM712_OUT));
      NOR2_X1 XNOR_3_3_NAND5_NUM712 (.ZN (XNOR_3_3_NAND5_NUM712_OUT), .A1 (XNOR_3_1_NAND5_NUM712_OUT), .A2 (XNOR_3_2_NAND5_NUM712_OUT));

      wire XNOR_4_1_NAND5_NUM712_OUT, XNOR_4_2_NAND5_NUM712_OUT, XNOR_4_3_NAND5_NUM712_OUT;
      NOR2_X1 XNOR_4_1_NAND5_NUM712 (.ZN (XNOR_4_1_NAND5_NUM712_OUT), .A1 (N1171), .A2 (GND));
      NOR2_X1 XNOR_4_2_NAND5_NUM712 (.ZN (XNOR_4_2_NAND5_NUM712_OUT), .A1 (GND), .A2 (XNOR_3_3_NAND5_NUM712_OUT));
      NOR2_X1 XNOR_4_3_NAND5_NUM712 (.ZN (XNOR_4_3_NAND5_NUM712_OUT), .A1 (XNOR_4_1_NAND5_NUM712_OUT), .A2 (XNOR_4_2_NAND5_NUM712_OUT));

      NOR2_X1 XNOR_5_1_NAND5_NUM712 (.ZN (N2543), .A1 (XNOR_4_3_NAND5_NUM712_OUT), .A2 (GND));
      wire XNOR_1_1_NAND5_NUM713_OUT, XNOR_1_2_NAND5_NUM713_OUT, XNOR_1_3_NAND5_NUM713_OUT;
      NOR2_X1 XNOR_1_1_NAND5_NUM713 (.ZN (XNOR_1_1_NAND5_NUM713_OUT), .A1 (N2286), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND5_NUM713 (.ZN (XNOR_1_2_NAND5_NUM713_OUT), .A1 (GND), .A2 (N2315));
      NOR2_X1 XNOR_1_3_NAND5_NUM713 (.ZN (XNOR_1_3_NAND5_NUM713_OUT), .A1 (XNOR_1_1_NAND5_NUM713_OUT), .A2 (XNOR_1_2_NAND5_NUM713_OUT));

      wire XNOR_2_1_NAND5_NUM713_OUT, XNOR_2_2_NAND5_NUM713_OUT, XNOR_2_3_NAND5_NUM713_OUT;
      NOR2_X1 XNOR_2_1_NAND5_NUM713 (.ZN (XNOR_2_1_NAND5_NUM713_OUT), .A1 (N2353), .A2 (GND));
      NOR2_X1 XNOR_2_2_NAND5_NUM713 (.ZN (XNOR_2_2_NAND5_NUM713_OUT), .A1 (GND), .A2 (N2104));
      NOR2_X1 XNOR_2_3_NAND5_NUM713 (.ZN (XNOR_2_3_NAND5_NUM713_OUT), .A1 (XNOR_2_1_NAND5_NUM713_OUT), .A2 (XNOR_2_2_NAND5_NUM713_OUT));

      wire XNOR_3_1_NAND5_NUM713_OUT, XNOR_3_2_NAND5_NUM713_OUT, XNOR_3_3_NAND5_NUM713_OUT;
      NOR2_X1 XNOR_3_1_NAND5_NUM713 (.ZN (XNOR_3_1_NAND5_NUM713_OUT), .A1 (XNOR_1_3_NAND5_NUM713_OUT), .A2 (GND));
      NOR2_X1 XNOR_3_2_NAND5_NUM713 (.ZN (XNOR_3_2_NAND5_NUM713_OUT), .A1 (GND), .A2 (XNOR_2_3_NAND5_NUM713_OUT));
      NOR2_X1 XNOR_3_3_NAND5_NUM713 (.ZN (XNOR_3_3_NAND5_NUM713_OUT), .A1 (XNOR_3_1_NAND5_NUM713_OUT), .A2 (XNOR_3_2_NAND5_NUM713_OUT));

      wire XNOR_4_1_NAND5_NUM713_OUT, XNOR_4_2_NAND5_NUM713_OUT, XNOR_4_3_NAND5_NUM713_OUT;
      NOR2_X1 XNOR_4_1_NAND5_NUM713 (.ZN (XNOR_4_1_NAND5_NUM713_OUT), .A1 (N1171), .A2 (GND));
      NOR2_X1 XNOR_4_2_NAND5_NUM713 (.ZN (XNOR_4_2_NAND5_NUM713_OUT), .A1 (GND), .A2 (XNOR_3_3_NAND5_NUM713_OUT));
      NOR2_X1 XNOR_4_3_NAND5_NUM713 (.ZN (XNOR_4_3_NAND5_NUM713_OUT), .A1 (XNOR_4_1_NAND5_NUM713_OUT), .A2 (XNOR_4_2_NAND5_NUM713_OUT));

      NOR2_X1 XNOR_5_1_NAND5_NUM713 (.ZN (N2546), .A1 (XNOR_4_3_NAND5_NUM713_OUT), .A2 (GND));
      wire XNOR_1_1_NAND5_NUM714_OUT, XNOR_1_2_NAND5_NUM714_OUT, XNOR_1_3_NAND5_NUM714_OUT;
      NOR2_X1 XNOR_1_1_NAND5_NUM714 (.ZN (XNOR_1_1_NAND5_NUM714_OUT), .A1 (N2297), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND5_NUM714 (.ZN (XNOR_1_2_NAND5_NUM714_OUT), .A1 (GND), .A2 (N2315));
      NOR2_X1 XNOR_1_3_NAND5_NUM714 (.ZN (XNOR_1_3_NAND5_NUM714_OUT), .A1 (XNOR_1_1_NAND5_NUM714_OUT), .A2 (XNOR_1_2_NAND5_NUM714_OUT));

      wire XNOR_2_1_NAND5_NUM714_OUT, XNOR_2_2_NAND5_NUM714_OUT, XNOR_2_3_NAND5_NUM714_OUT;
      NOR2_X1 XNOR_2_1_NAND5_NUM714 (.ZN (XNOR_2_1_NAND5_NUM714_OUT), .A1 (N2375), .A2 (GND));
      NOR2_X1 XNOR_2_2_NAND5_NUM714 (.ZN (XNOR_2_2_NAND5_NUM714_OUT), .A1 (GND), .A2 (N2119));
      NOR2_X1 XNOR_2_3_NAND5_NUM714 (.ZN (XNOR_2_3_NAND5_NUM714_OUT), .A1 (XNOR_2_1_NAND5_NUM714_OUT), .A2 (XNOR_2_2_NAND5_NUM714_OUT));

      wire XNOR_3_1_NAND5_NUM714_OUT, XNOR_3_2_NAND5_NUM714_OUT, XNOR_3_3_NAND5_NUM714_OUT;
      NOR2_X1 XNOR_3_1_NAND5_NUM714 (.ZN (XNOR_3_1_NAND5_NUM714_OUT), .A1 (XNOR_1_3_NAND5_NUM714_OUT), .A2 (GND));
      NOR2_X1 XNOR_3_2_NAND5_NUM714 (.ZN (XNOR_3_2_NAND5_NUM714_OUT), .A1 (GND), .A2 (XNOR_2_3_NAND5_NUM714_OUT));
      NOR2_X1 XNOR_3_3_NAND5_NUM714 (.ZN (XNOR_3_3_NAND5_NUM714_OUT), .A1 (XNOR_3_1_NAND5_NUM714_OUT), .A2 (XNOR_3_2_NAND5_NUM714_OUT));

      wire XNOR_4_1_NAND5_NUM714_OUT, XNOR_4_2_NAND5_NUM714_OUT, XNOR_4_3_NAND5_NUM714_OUT;
      NOR2_X1 XNOR_4_1_NAND5_NUM714 (.ZN (XNOR_4_1_NAND5_NUM714_OUT), .A1 (N1188), .A2 (GND));
      NOR2_X1 XNOR_4_2_NAND5_NUM714 (.ZN (XNOR_4_2_NAND5_NUM714_OUT), .A1 (GND), .A2 (XNOR_3_3_NAND5_NUM714_OUT));
      NOR2_X1 XNOR_4_3_NAND5_NUM714 (.ZN (XNOR_4_3_NAND5_NUM714_OUT), .A1 (XNOR_4_1_NAND5_NUM714_OUT), .A2 (XNOR_4_2_NAND5_NUM714_OUT));

      NOR2_X1 XNOR_5_1_NAND5_NUM714 (.ZN (N2549), .A1 (XNOR_4_3_NAND5_NUM714_OUT), .A2 (GND));
      wire XNOR_1_1_NAND5_NUM715_OUT, XNOR_1_2_NAND5_NUM715_OUT, XNOR_1_3_NAND5_NUM715_OUT;
      NOR2_X1 XNOR_1_1_NAND5_NUM715 (.ZN (XNOR_1_1_NAND5_NUM715_OUT), .A1 (N2297), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND5_NUM715 (.ZN (XNOR_1_2_NAND5_NUM715_OUT), .A1 (GND), .A2 (N2326));
      NOR2_X1 XNOR_1_3_NAND5_NUM715 (.ZN (XNOR_1_3_NAND5_NUM715_OUT), .A1 (XNOR_1_1_NAND5_NUM715_OUT), .A2 (XNOR_1_2_NAND5_NUM715_OUT));

      wire XNOR_2_1_NAND5_NUM715_OUT, XNOR_2_2_NAND5_NUM715_OUT, XNOR_2_3_NAND5_NUM715_OUT;
      NOR2_X1 XNOR_2_1_NAND5_NUM715 (.ZN (XNOR_2_1_NAND5_NUM715_OUT), .A1 (N2361), .A2 (GND));
      NOR2_X1 XNOR_2_2_NAND5_NUM715 (.ZN (XNOR_2_2_NAND5_NUM715_OUT), .A1 (GND), .A2 (N2143));
      NOR2_X1 XNOR_2_3_NAND5_NUM715 (.ZN (XNOR_2_3_NAND5_NUM715_OUT), .A1 (XNOR_2_1_NAND5_NUM715_OUT), .A2 (XNOR_2_2_NAND5_NUM715_OUT));

      wire XNOR_3_1_NAND5_NUM715_OUT, XNOR_3_2_NAND5_NUM715_OUT, XNOR_3_3_NAND5_NUM715_OUT;
      NOR2_X1 XNOR_3_1_NAND5_NUM715 (.ZN (XNOR_3_1_NAND5_NUM715_OUT), .A1 (XNOR_1_3_NAND5_NUM715_OUT), .A2 (GND));
      NOR2_X1 XNOR_3_2_NAND5_NUM715 (.ZN (XNOR_3_2_NAND5_NUM715_OUT), .A1 (GND), .A2 (XNOR_2_3_NAND5_NUM715_OUT));
      NOR2_X1 XNOR_3_3_NAND5_NUM715 (.ZN (XNOR_3_3_NAND5_NUM715_OUT), .A1 (XNOR_3_1_NAND5_NUM715_OUT), .A2 (XNOR_3_2_NAND5_NUM715_OUT));

      wire XNOR_4_1_NAND5_NUM715_OUT, XNOR_4_2_NAND5_NUM715_OUT, XNOR_4_3_NAND5_NUM715_OUT;
      NOR2_X1 XNOR_4_1_NAND5_NUM715 (.ZN (XNOR_4_1_NAND5_NUM715_OUT), .A1 (N1188), .A2 (GND));
      NOR2_X1 XNOR_4_2_NAND5_NUM715 (.ZN (XNOR_4_2_NAND5_NUM715_OUT), .A1 (GND), .A2 (XNOR_3_3_NAND5_NUM715_OUT));
      NOR2_X1 XNOR_4_3_NAND5_NUM715 (.ZN (XNOR_4_3_NAND5_NUM715_OUT), .A1 (XNOR_4_1_NAND5_NUM715_OUT), .A2 (XNOR_4_2_NAND5_NUM715_OUT));

      NOR2_X1 XNOR_5_1_NAND5_NUM715 (.ZN (N2552), .A1 (XNOR_4_3_NAND5_NUM715_OUT), .A2 (GND));
      wire XNOR_1_1_NAND5_NUM716_OUT, XNOR_1_2_NAND5_NUM716_OUT, XNOR_1_3_NAND5_NUM716_OUT;
      NOR2_X1 XNOR_1_1_NAND5_NUM716 (.ZN (XNOR_1_1_NAND5_NUM716_OUT), .A1 (N2297), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND5_NUM716 (.ZN (XNOR_1_2_NAND5_NUM716_OUT), .A1 (GND), .A2 (N2326));
      NOR2_X1 XNOR_1_3_NAND5_NUM716 (.ZN (XNOR_1_3_NAND5_NUM716_OUT), .A1 (XNOR_1_1_NAND5_NUM716_OUT), .A2 (XNOR_1_2_NAND5_NUM716_OUT));

      wire XNOR_2_1_NAND5_NUM716_OUT, XNOR_2_2_NAND5_NUM716_OUT, XNOR_2_3_NAND5_NUM716_OUT;
      NOR2_X1 XNOR_2_1_NAND5_NUM716 (.ZN (XNOR_2_1_NAND5_NUM716_OUT), .A1 (N2375), .A2 (GND));
      NOR2_X1 XNOR_2_2_NAND5_NUM716 (.ZN (XNOR_2_2_NAND5_NUM716_OUT), .A1 (GND), .A2 (N2129));
      NOR2_X1 XNOR_2_3_NAND5_NUM716 (.ZN (XNOR_2_3_NAND5_NUM716_OUT), .A1 (XNOR_2_1_NAND5_NUM716_OUT), .A2 (XNOR_2_2_NAND5_NUM716_OUT));

      wire XNOR_3_1_NAND5_NUM716_OUT, XNOR_3_2_NAND5_NUM716_OUT, XNOR_3_3_NAND5_NUM716_OUT;
      NOR2_X1 XNOR_3_1_NAND5_NUM716 (.ZN (XNOR_3_1_NAND5_NUM716_OUT), .A1 (XNOR_1_3_NAND5_NUM716_OUT), .A2 (GND));
      NOR2_X1 XNOR_3_2_NAND5_NUM716 (.ZN (XNOR_3_2_NAND5_NUM716_OUT), .A1 (GND), .A2 (XNOR_2_3_NAND5_NUM716_OUT));
      NOR2_X1 XNOR_3_3_NAND5_NUM716 (.ZN (XNOR_3_3_NAND5_NUM716_OUT), .A1 (XNOR_3_1_NAND5_NUM716_OUT), .A2 (XNOR_3_2_NAND5_NUM716_OUT));

      wire XNOR_4_1_NAND5_NUM716_OUT, XNOR_4_2_NAND5_NUM716_OUT, XNOR_4_3_NAND5_NUM716_OUT;
      NOR2_X1 XNOR_4_1_NAND5_NUM716 (.ZN (XNOR_4_1_NAND5_NUM716_OUT), .A1 (N1188), .A2 (GND));
      NOR2_X1 XNOR_4_2_NAND5_NUM716 (.ZN (XNOR_4_2_NAND5_NUM716_OUT), .A1 (GND), .A2 (XNOR_3_3_NAND5_NUM716_OUT));
      NOR2_X1 XNOR_4_3_NAND5_NUM716 (.ZN (XNOR_4_3_NAND5_NUM716_OUT), .A1 (XNOR_4_1_NAND5_NUM716_OUT), .A2 (XNOR_4_2_NAND5_NUM716_OUT));

      NOR2_X1 XNOR_5_1_NAND5_NUM716 (.ZN (N2555), .A1 (XNOR_4_3_NAND5_NUM716_OUT), .A2 (GND));
      wire XNOR_1_1_AND5_NUM717_OUT, XNOR_1_2_AND5_NUM717_OUT, XNOR_1_3_AND5_NUM717_OUT;
      NOR2_X1 XNOR_1_1_AND5_NUM717 (.ZN (XNOR_1_1_AND5_NUM717_OUT), .A1 (N2286), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND5_NUM717 (.ZN (XNOR_1_2_AND5_NUM717_OUT), .A1 (GND), .A2 (N2315));
      NOR2_X1 XNOR_1_3_AND5_NUM717 (.ZN (XNOR_1_3_AND5_NUM717_OUT), .A1 (XNOR_1_1_AND5_NUM717_OUT), .A2 (XNOR_1_2_AND5_NUM717_OUT));

      wire XNOR_2_1_AND5_NUM717_OUT, XNOR_2_2_AND5_NUM717_OUT, XNOR_2_3_AND5_NUM717_OUT;
      NOR2_X1 XNOR_2_1_AND5_NUM717 (.ZN (XNOR_2_1_AND5_NUM717_OUT), .A1 (N2361), .A2 (GND));
      NOR2_X1 XNOR_2_2_AND5_NUM717 (.ZN (XNOR_2_2_AND5_NUM717_OUT), .A1 (GND), .A2 (N2104));
      NOR2_X1 XNOR_2_3_AND5_NUM717 (.ZN (XNOR_2_3_AND5_NUM717_OUT), .A1 (XNOR_2_1_AND5_NUM717_OUT), .A2 (XNOR_2_2_AND5_NUM717_OUT));

      wire XNOR_3_1_AND5_NUM717_OUT, XNOR_3_2_AND5_NUM717_OUT, XNOR_3_3_AND5_NUM717_OUT;
      NOR2_X1 XNOR_3_1_AND5_NUM717 (.ZN (XNOR_3_1_AND5_NUM717_OUT), .A1 (XNOR_1_3_AND5_NUM717_OUT), .A2 (GND));
      NOR2_X1 XNOR_3_2_AND5_NUM717 (.ZN (XNOR_3_2_AND5_NUM717_OUT), .A1 (GND), .A2 (XNOR_2_3_AND5_NUM717_OUT));
      NOR2_X1 XNOR_3_3_AND5_NUM717 (.ZN (XNOR_3_3_AND5_NUM717_OUT), .A1 (XNOR_3_1_AND5_NUM717_OUT), .A2 (XNOR_3_2_AND5_NUM717_OUT));

      wire XNOR_4_1_AND5_NUM717_OUT, XNOR_4_2_AND5_NUM717_OUT;
      NOR2_X1 XNOR_4_1_AND5_NUM717 (.ZN (XNOR_4_1_AND5_NUM717_OUT), .A1 (N1171), .A2 (GND));
      NOR2_X1 XNOR_4_2_AND5_NUM717 (.ZN (XNOR_4_2_AND5_NUM717_OUT), .A1 (GND), .A2 (XNOR_3_3_AND5_NUM717_OUT));
      NOR2_X1 XNOR_4_3_AND5_NUM717 (.ZN (N2558), .A1 (XNOR_4_1_AND5_NUM717_OUT), .A2 (XNOR_4_2_AND5_NUM717_OUT));
      wire XNOR_1_1_AND5_NUM718_OUT, XNOR_1_2_AND5_NUM718_OUT, XNOR_1_3_AND5_NUM718_OUT;
      NOR2_X1 XNOR_1_1_AND5_NUM718 (.ZN (XNOR_1_1_AND5_NUM718_OUT), .A1 (N2286), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND5_NUM718 (.ZN (XNOR_1_2_AND5_NUM718_OUT), .A1 (GND), .A2 (N2315));
      NOR2_X1 XNOR_1_3_AND5_NUM718 (.ZN (XNOR_1_3_AND5_NUM718_OUT), .A1 (XNOR_1_1_AND5_NUM718_OUT), .A2 (XNOR_1_2_AND5_NUM718_OUT));

      wire XNOR_2_1_AND5_NUM718_OUT, XNOR_2_2_AND5_NUM718_OUT, XNOR_2_3_AND5_NUM718_OUT;
      NOR2_X1 XNOR_2_1_AND5_NUM718 (.ZN (XNOR_2_1_AND5_NUM718_OUT), .A1 (N2340), .A2 (GND));
      NOR2_X1 XNOR_2_2_AND5_NUM718 (.ZN (XNOR_2_2_AND5_NUM718_OUT), .A1 (GND), .A2 (N2129));
      NOR2_X1 XNOR_2_3_AND5_NUM718 (.ZN (XNOR_2_3_AND5_NUM718_OUT), .A1 (XNOR_2_1_AND5_NUM718_OUT), .A2 (XNOR_2_2_AND5_NUM718_OUT));

      wire XNOR_3_1_AND5_NUM718_OUT, XNOR_3_2_AND5_NUM718_OUT, XNOR_3_3_AND5_NUM718_OUT;
      NOR2_X1 XNOR_3_1_AND5_NUM718 (.ZN (XNOR_3_1_AND5_NUM718_OUT), .A1 (XNOR_1_3_AND5_NUM718_OUT), .A2 (GND));
      NOR2_X1 XNOR_3_2_AND5_NUM718 (.ZN (XNOR_3_2_AND5_NUM718_OUT), .A1 (GND), .A2 (XNOR_2_3_AND5_NUM718_OUT));
      NOR2_X1 XNOR_3_3_AND5_NUM718 (.ZN (XNOR_3_3_AND5_NUM718_OUT), .A1 (XNOR_3_1_AND5_NUM718_OUT), .A2 (XNOR_3_2_AND5_NUM718_OUT));

      wire XNOR_4_1_AND5_NUM718_OUT, XNOR_4_2_AND5_NUM718_OUT;
      NOR2_X1 XNOR_4_1_AND5_NUM718 (.ZN (XNOR_4_1_AND5_NUM718_OUT), .A1 (N1171), .A2 (GND));
      NOR2_X1 XNOR_4_2_AND5_NUM718 (.ZN (XNOR_4_2_AND5_NUM718_OUT), .A1 (GND), .A2 (XNOR_3_3_AND5_NUM718_OUT));
      NOR2_X1 XNOR_4_3_AND5_NUM718 (.ZN (N2561), .A1 (XNOR_4_1_AND5_NUM718_OUT), .A2 (XNOR_4_2_AND5_NUM718_OUT));
      wire XNOR_1_1_AND5_NUM719_OUT, XNOR_1_2_AND5_NUM719_OUT, XNOR_1_3_AND5_NUM719_OUT;
      NOR2_X1 XNOR_1_1_AND5_NUM719 (.ZN (XNOR_1_1_AND5_NUM719_OUT), .A1 (N2286), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND5_NUM719 (.ZN (XNOR_1_2_AND5_NUM719_OUT), .A1 (GND), .A2 (N2315));
      NOR2_X1 XNOR_1_3_AND5_NUM719 (.ZN (XNOR_1_3_AND5_NUM719_OUT), .A1 (XNOR_1_1_AND5_NUM719_OUT), .A2 (XNOR_1_2_AND5_NUM719_OUT));

      wire XNOR_2_1_AND5_NUM719_OUT, XNOR_2_2_AND5_NUM719_OUT, XNOR_2_3_AND5_NUM719_OUT;
      NOR2_X1 XNOR_2_1_AND5_NUM719 (.ZN (XNOR_2_1_AND5_NUM719_OUT), .A1 (N2340), .A2 (GND));
      NOR2_X1 XNOR_2_2_AND5_NUM719 (.ZN (XNOR_2_2_AND5_NUM719_OUT), .A1 (GND), .A2 (N2119));
      NOR2_X1 XNOR_2_3_AND5_NUM719 (.ZN (XNOR_2_3_AND5_NUM719_OUT), .A1 (XNOR_2_1_AND5_NUM719_OUT), .A2 (XNOR_2_2_AND5_NUM719_OUT));

      wire XNOR_3_1_AND5_NUM719_OUT, XNOR_3_2_AND5_NUM719_OUT, XNOR_3_3_AND5_NUM719_OUT;
      NOR2_X1 XNOR_3_1_AND5_NUM719 (.ZN (XNOR_3_1_AND5_NUM719_OUT), .A1 (XNOR_1_3_AND5_NUM719_OUT), .A2 (GND));
      NOR2_X1 XNOR_3_2_AND5_NUM719 (.ZN (XNOR_3_2_AND5_NUM719_OUT), .A1 (GND), .A2 (XNOR_2_3_AND5_NUM719_OUT));
      NOR2_X1 XNOR_3_3_AND5_NUM719 (.ZN (XNOR_3_3_AND5_NUM719_OUT), .A1 (XNOR_3_1_AND5_NUM719_OUT), .A2 (XNOR_3_2_AND5_NUM719_OUT));

      wire XNOR_4_1_AND5_NUM719_OUT, XNOR_4_2_AND5_NUM719_OUT;
      NOR2_X1 XNOR_4_1_AND5_NUM719 (.ZN (XNOR_4_1_AND5_NUM719_OUT), .A1 (N1171), .A2 (GND));
      NOR2_X1 XNOR_4_2_AND5_NUM719 (.ZN (XNOR_4_2_AND5_NUM719_OUT), .A1 (GND), .A2 (XNOR_3_3_AND5_NUM719_OUT));
      NOR2_X1 XNOR_4_3_AND5_NUM719 (.ZN (N2564), .A1 (XNOR_4_1_AND5_NUM719_OUT), .A2 (XNOR_4_2_AND5_NUM719_OUT));
      wire XNOR_1_1_AND5_NUM720_OUT, XNOR_1_2_AND5_NUM720_OUT, XNOR_1_3_AND5_NUM720_OUT;
      NOR2_X1 XNOR_1_1_AND5_NUM720 (.ZN (XNOR_1_1_AND5_NUM720_OUT), .A1 (N2286), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND5_NUM720 (.ZN (XNOR_1_2_AND5_NUM720_OUT), .A1 (GND), .A2 (N2315));
      NOR2_X1 XNOR_1_3_AND5_NUM720 (.ZN (XNOR_1_3_AND5_NUM720_OUT), .A1 (XNOR_1_1_AND5_NUM720_OUT), .A2 (XNOR_1_2_AND5_NUM720_OUT));

      wire XNOR_2_1_AND5_NUM720_OUT, XNOR_2_2_AND5_NUM720_OUT, XNOR_2_3_AND5_NUM720_OUT;
      NOR2_X1 XNOR_2_1_AND5_NUM720 (.ZN (XNOR_2_1_AND5_NUM720_OUT), .A1 (N2353), .A2 (GND));
      NOR2_X1 XNOR_2_2_AND5_NUM720 (.ZN (XNOR_2_2_AND5_NUM720_OUT), .A1 (GND), .A2 (N2104));
      NOR2_X1 XNOR_2_3_AND5_NUM720 (.ZN (XNOR_2_3_AND5_NUM720_OUT), .A1 (XNOR_2_1_AND5_NUM720_OUT), .A2 (XNOR_2_2_AND5_NUM720_OUT));

      wire XNOR_3_1_AND5_NUM720_OUT, XNOR_3_2_AND5_NUM720_OUT, XNOR_3_3_AND5_NUM720_OUT;
      NOR2_X1 XNOR_3_1_AND5_NUM720 (.ZN (XNOR_3_1_AND5_NUM720_OUT), .A1 (XNOR_1_3_AND5_NUM720_OUT), .A2 (GND));
      NOR2_X1 XNOR_3_2_AND5_NUM720 (.ZN (XNOR_3_2_AND5_NUM720_OUT), .A1 (GND), .A2 (XNOR_2_3_AND5_NUM720_OUT));
      NOR2_X1 XNOR_3_3_AND5_NUM720 (.ZN (XNOR_3_3_AND5_NUM720_OUT), .A1 (XNOR_3_1_AND5_NUM720_OUT), .A2 (XNOR_3_2_AND5_NUM720_OUT));

      wire XNOR_4_1_AND5_NUM720_OUT, XNOR_4_2_AND5_NUM720_OUT;
      NOR2_X1 XNOR_4_1_AND5_NUM720 (.ZN (XNOR_4_1_AND5_NUM720_OUT), .A1 (N1171), .A2 (GND));
      NOR2_X1 XNOR_4_2_AND5_NUM720 (.ZN (XNOR_4_2_AND5_NUM720_OUT), .A1 (GND), .A2 (XNOR_3_3_AND5_NUM720_OUT));
      NOR2_X1 XNOR_4_3_AND5_NUM720 (.ZN (N2567), .A1 (XNOR_4_1_AND5_NUM720_OUT), .A2 (XNOR_4_2_AND5_NUM720_OUT));
      wire XNOR_1_1_AND5_NUM721_OUT, XNOR_1_2_AND5_NUM721_OUT, XNOR_1_3_AND5_NUM721_OUT;
      NOR2_X1 XNOR_1_1_AND5_NUM721 (.ZN (XNOR_1_1_AND5_NUM721_OUT), .A1 (N2297), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND5_NUM721 (.ZN (XNOR_1_2_AND5_NUM721_OUT), .A1 (GND), .A2 (N2315));
      NOR2_X1 XNOR_1_3_AND5_NUM721 (.ZN (XNOR_1_3_AND5_NUM721_OUT), .A1 (XNOR_1_1_AND5_NUM721_OUT), .A2 (XNOR_1_2_AND5_NUM721_OUT));

      wire XNOR_2_1_AND5_NUM721_OUT, XNOR_2_2_AND5_NUM721_OUT, XNOR_2_3_AND5_NUM721_OUT;
      NOR2_X1 XNOR_2_1_AND5_NUM721 (.ZN (XNOR_2_1_AND5_NUM721_OUT), .A1 (N2375), .A2 (GND));
      NOR2_X1 XNOR_2_2_AND5_NUM721 (.ZN (XNOR_2_2_AND5_NUM721_OUT), .A1 (GND), .A2 (N2119));
      NOR2_X1 XNOR_2_3_AND5_NUM721 (.ZN (XNOR_2_3_AND5_NUM721_OUT), .A1 (XNOR_2_1_AND5_NUM721_OUT), .A2 (XNOR_2_2_AND5_NUM721_OUT));

      wire XNOR_3_1_AND5_NUM721_OUT, XNOR_3_2_AND5_NUM721_OUT, XNOR_3_3_AND5_NUM721_OUT;
      NOR2_X1 XNOR_3_1_AND5_NUM721 (.ZN (XNOR_3_1_AND5_NUM721_OUT), .A1 (XNOR_1_3_AND5_NUM721_OUT), .A2 (GND));
      NOR2_X1 XNOR_3_2_AND5_NUM721 (.ZN (XNOR_3_2_AND5_NUM721_OUT), .A1 (GND), .A2 (XNOR_2_3_AND5_NUM721_OUT));
      NOR2_X1 XNOR_3_3_AND5_NUM721 (.ZN (XNOR_3_3_AND5_NUM721_OUT), .A1 (XNOR_3_1_AND5_NUM721_OUT), .A2 (XNOR_3_2_AND5_NUM721_OUT));

      wire XNOR_4_1_AND5_NUM721_OUT, XNOR_4_2_AND5_NUM721_OUT;
      NOR2_X1 XNOR_4_1_AND5_NUM721 (.ZN (XNOR_4_1_AND5_NUM721_OUT), .A1 (N1188), .A2 (GND));
      NOR2_X1 XNOR_4_2_AND5_NUM721 (.ZN (XNOR_4_2_AND5_NUM721_OUT), .A1 (GND), .A2 (XNOR_3_3_AND5_NUM721_OUT));
      NOR2_X1 XNOR_4_3_AND5_NUM721 (.ZN (N2570), .A1 (XNOR_4_1_AND5_NUM721_OUT), .A2 (XNOR_4_2_AND5_NUM721_OUT));
      wire XNOR_1_1_AND5_NUM722_OUT, XNOR_1_2_AND5_NUM722_OUT, XNOR_1_3_AND5_NUM722_OUT;
      NOR2_X1 XNOR_1_1_AND5_NUM722 (.ZN (XNOR_1_1_AND5_NUM722_OUT), .A1 (N2297), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND5_NUM722 (.ZN (XNOR_1_2_AND5_NUM722_OUT), .A1 (GND), .A2 (N2326));
      NOR2_X1 XNOR_1_3_AND5_NUM722 (.ZN (XNOR_1_3_AND5_NUM722_OUT), .A1 (XNOR_1_1_AND5_NUM722_OUT), .A2 (XNOR_1_2_AND5_NUM722_OUT));

      wire XNOR_2_1_AND5_NUM722_OUT, XNOR_2_2_AND5_NUM722_OUT, XNOR_2_3_AND5_NUM722_OUT;
      NOR2_X1 XNOR_2_1_AND5_NUM722 (.ZN (XNOR_2_1_AND5_NUM722_OUT), .A1 (N2361), .A2 (GND));
      NOR2_X1 XNOR_2_2_AND5_NUM722 (.ZN (XNOR_2_2_AND5_NUM722_OUT), .A1 (GND), .A2 (N2143));
      NOR2_X1 XNOR_2_3_AND5_NUM722 (.ZN (XNOR_2_3_AND5_NUM722_OUT), .A1 (XNOR_2_1_AND5_NUM722_OUT), .A2 (XNOR_2_2_AND5_NUM722_OUT));

      wire XNOR_3_1_AND5_NUM722_OUT, XNOR_3_2_AND5_NUM722_OUT, XNOR_3_3_AND5_NUM722_OUT;
      NOR2_X1 XNOR_3_1_AND5_NUM722 (.ZN (XNOR_3_1_AND5_NUM722_OUT), .A1 (XNOR_1_3_AND5_NUM722_OUT), .A2 (GND));
      NOR2_X1 XNOR_3_2_AND5_NUM722 (.ZN (XNOR_3_2_AND5_NUM722_OUT), .A1 (GND), .A2 (XNOR_2_3_AND5_NUM722_OUT));
      NOR2_X1 XNOR_3_3_AND5_NUM722 (.ZN (XNOR_3_3_AND5_NUM722_OUT), .A1 (XNOR_3_1_AND5_NUM722_OUT), .A2 (XNOR_3_2_AND5_NUM722_OUT));

      wire XNOR_4_1_AND5_NUM722_OUT, XNOR_4_2_AND5_NUM722_OUT;
      NOR2_X1 XNOR_4_1_AND5_NUM722 (.ZN (XNOR_4_1_AND5_NUM722_OUT), .A1 (N1188), .A2 (GND));
      NOR2_X1 XNOR_4_2_AND5_NUM722 (.ZN (XNOR_4_2_AND5_NUM722_OUT), .A1 (GND), .A2 (XNOR_3_3_AND5_NUM722_OUT));
      NOR2_X1 XNOR_4_3_AND5_NUM722 (.ZN (N2573), .A1 (XNOR_4_1_AND5_NUM722_OUT), .A2 (XNOR_4_2_AND5_NUM722_OUT));
      wire XNOR_1_1_AND5_NUM723_OUT, XNOR_1_2_AND5_NUM723_OUT, XNOR_1_3_AND5_NUM723_OUT;
      NOR2_X1 XNOR_1_1_AND5_NUM723 (.ZN (XNOR_1_1_AND5_NUM723_OUT), .A1 (N2297), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND5_NUM723 (.ZN (XNOR_1_2_AND5_NUM723_OUT), .A1 (GND), .A2 (N2326));
      NOR2_X1 XNOR_1_3_AND5_NUM723 (.ZN (XNOR_1_3_AND5_NUM723_OUT), .A1 (XNOR_1_1_AND5_NUM723_OUT), .A2 (XNOR_1_2_AND5_NUM723_OUT));

      wire XNOR_2_1_AND5_NUM723_OUT, XNOR_2_2_AND5_NUM723_OUT, XNOR_2_3_AND5_NUM723_OUT;
      NOR2_X1 XNOR_2_1_AND5_NUM723 (.ZN (XNOR_2_1_AND5_NUM723_OUT), .A1 (N2375), .A2 (GND));
      NOR2_X1 XNOR_2_2_AND5_NUM723 (.ZN (XNOR_2_2_AND5_NUM723_OUT), .A1 (GND), .A2 (N2129));
      NOR2_X1 XNOR_2_3_AND5_NUM723 (.ZN (XNOR_2_3_AND5_NUM723_OUT), .A1 (XNOR_2_1_AND5_NUM723_OUT), .A2 (XNOR_2_2_AND5_NUM723_OUT));

      wire XNOR_3_1_AND5_NUM723_OUT, XNOR_3_2_AND5_NUM723_OUT, XNOR_3_3_AND5_NUM723_OUT;
      NOR2_X1 XNOR_3_1_AND5_NUM723 (.ZN (XNOR_3_1_AND5_NUM723_OUT), .A1 (XNOR_1_3_AND5_NUM723_OUT), .A2 (GND));
      NOR2_X1 XNOR_3_2_AND5_NUM723 (.ZN (XNOR_3_2_AND5_NUM723_OUT), .A1 (GND), .A2 (XNOR_2_3_AND5_NUM723_OUT));
      NOR2_X1 XNOR_3_3_AND5_NUM723 (.ZN (XNOR_3_3_AND5_NUM723_OUT), .A1 (XNOR_3_1_AND5_NUM723_OUT), .A2 (XNOR_3_2_AND5_NUM723_OUT));

      wire XNOR_4_1_AND5_NUM723_OUT, XNOR_4_2_AND5_NUM723_OUT;
      NOR2_X1 XNOR_4_1_AND5_NUM723 (.ZN (XNOR_4_1_AND5_NUM723_OUT), .A1 (N1188), .A2 (GND));
      NOR2_X1 XNOR_4_2_AND5_NUM723 (.ZN (XNOR_4_2_AND5_NUM723_OUT), .A1 (GND), .A2 (XNOR_3_3_AND5_NUM723_OUT));
      NOR2_X1 XNOR_4_3_AND5_NUM723 (.ZN (N2576), .A1 (XNOR_4_1_AND5_NUM723_OUT), .A2 (XNOR_4_2_AND5_NUM723_OUT));
      wire XNOR_1_1_NAND5_NUM724_OUT, XNOR_1_2_NAND5_NUM724_OUT, XNOR_1_3_NAND5_NUM724_OUT;
      NOR2_X1 XNOR_1_1_NAND5_NUM724 (.ZN (XNOR_1_1_NAND5_NUM724_OUT), .A1 (N2286), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND5_NUM724 (.ZN (XNOR_1_2_NAND5_NUM724_OUT), .A1 (GND), .A2 (N2427));
      NOR2_X1 XNOR_1_3_NAND5_NUM724 (.ZN (XNOR_1_3_NAND5_NUM724_OUT), .A1 (XNOR_1_1_NAND5_NUM724_OUT), .A2 (XNOR_1_2_NAND5_NUM724_OUT));

      wire XNOR_2_1_NAND5_NUM724_OUT, XNOR_2_2_NAND5_NUM724_OUT, XNOR_2_3_NAND5_NUM724_OUT;
      NOR2_X1 XNOR_2_1_NAND5_NUM724 (.ZN (XNOR_2_1_NAND5_NUM724_OUT), .A1 (N2361), .A2 (GND));
      NOR2_X1 XNOR_2_2_NAND5_NUM724 (.ZN (XNOR_2_2_NAND5_NUM724_OUT), .A1 (GND), .A2 (N2129));
      NOR2_X1 XNOR_2_3_NAND5_NUM724 (.ZN (XNOR_2_3_NAND5_NUM724_OUT), .A1 (XNOR_2_1_NAND5_NUM724_OUT), .A2 (XNOR_2_2_NAND5_NUM724_OUT));

      wire XNOR_3_1_NAND5_NUM724_OUT, XNOR_3_2_NAND5_NUM724_OUT, XNOR_3_3_NAND5_NUM724_OUT;
      NOR2_X1 XNOR_3_1_NAND5_NUM724 (.ZN (XNOR_3_1_NAND5_NUM724_OUT), .A1 (XNOR_1_3_NAND5_NUM724_OUT), .A2 (GND));
      NOR2_X1 XNOR_3_2_NAND5_NUM724 (.ZN (XNOR_3_2_NAND5_NUM724_OUT), .A1 (GND), .A2 (XNOR_2_3_NAND5_NUM724_OUT));
      NOR2_X1 XNOR_3_3_NAND5_NUM724 (.ZN (XNOR_3_3_NAND5_NUM724_OUT), .A1 (XNOR_3_1_NAND5_NUM724_OUT), .A2 (XNOR_3_2_NAND5_NUM724_OUT));

      wire XNOR_4_1_NAND5_NUM724_OUT, XNOR_4_2_NAND5_NUM724_OUT, XNOR_4_3_NAND5_NUM724_OUT;
      NOR2_X1 XNOR_4_1_NAND5_NUM724 (.ZN (XNOR_4_1_NAND5_NUM724_OUT), .A1 (N1171), .A2 (GND));
      NOR2_X1 XNOR_4_2_NAND5_NUM724 (.ZN (XNOR_4_2_NAND5_NUM724_OUT), .A1 (GND), .A2 (XNOR_3_3_NAND5_NUM724_OUT));
      NOR2_X1 XNOR_4_3_NAND5_NUM724 (.ZN (XNOR_4_3_NAND5_NUM724_OUT), .A1 (XNOR_4_1_NAND5_NUM724_OUT), .A2 (XNOR_4_2_NAND5_NUM724_OUT));

      NOR2_X1 XNOR_5_1_NAND5_NUM724 (.ZN (N2594), .A1 (XNOR_4_3_NAND5_NUM724_OUT), .A2 (GND));
      wire XNOR_1_1_NAND5_NUM725_OUT, XNOR_1_2_NAND5_NUM725_OUT, XNOR_1_3_NAND5_NUM725_OUT;
      NOR2_X1 XNOR_1_1_NAND5_NUM725 (.ZN (XNOR_1_1_NAND5_NUM725_OUT), .A1 (N2297), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND5_NUM725 (.ZN (XNOR_1_2_NAND5_NUM725_OUT), .A1 (GND), .A2 (N2427));
      NOR2_X1 XNOR_1_3_NAND5_NUM725 (.ZN (XNOR_1_3_NAND5_NUM725_OUT), .A1 (XNOR_1_1_NAND5_NUM725_OUT), .A2 (XNOR_1_2_NAND5_NUM725_OUT));

      wire XNOR_2_1_NAND5_NUM725_OUT, XNOR_2_2_NAND5_NUM725_OUT, XNOR_2_3_NAND5_NUM725_OUT;
      NOR2_X1 XNOR_2_1_NAND5_NUM725 (.ZN (XNOR_2_1_NAND5_NUM725_OUT), .A1 (N2361), .A2 (GND));
      NOR2_X1 XNOR_2_2_NAND5_NUM725 (.ZN (XNOR_2_2_NAND5_NUM725_OUT), .A1 (GND), .A2 (N2119));
      NOR2_X1 XNOR_2_3_NAND5_NUM725 (.ZN (XNOR_2_3_NAND5_NUM725_OUT), .A1 (XNOR_2_1_NAND5_NUM725_OUT), .A2 (XNOR_2_2_NAND5_NUM725_OUT));

      wire XNOR_3_1_NAND5_NUM725_OUT, XNOR_3_2_NAND5_NUM725_OUT, XNOR_3_3_NAND5_NUM725_OUT;
      NOR2_X1 XNOR_3_1_NAND5_NUM725 (.ZN (XNOR_3_1_NAND5_NUM725_OUT), .A1 (XNOR_1_3_NAND5_NUM725_OUT), .A2 (GND));
      NOR2_X1 XNOR_3_2_NAND5_NUM725 (.ZN (XNOR_3_2_NAND5_NUM725_OUT), .A1 (GND), .A2 (XNOR_2_3_NAND5_NUM725_OUT));
      NOR2_X1 XNOR_3_3_NAND5_NUM725 (.ZN (XNOR_3_3_NAND5_NUM725_OUT), .A1 (XNOR_3_1_NAND5_NUM725_OUT), .A2 (XNOR_3_2_NAND5_NUM725_OUT));

      wire XNOR_4_1_NAND5_NUM725_OUT, XNOR_4_2_NAND5_NUM725_OUT, XNOR_4_3_NAND5_NUM725_OUT;
      NOR2_X1 XNOR_4_1_NAND5_NUM725 (.ZN (XNOR_4_1_NAND5_NUM725_OUT), .A1 (N1171), .A2 (GND));
      NOR2_X1 XNOR_4_2_NAND5_NUM725 (.ZN (XNOR_4_2_NAND5_NUM725_OUT), .A1 (GND), .A2 (XNOR_3_3_NAND5_NUM725_OUT));
      NOR2_X1 XNOR_4_3_NAND5_NUM725 (.ZN (XNOR_4_3_NAND5_NUM725_OUT), .A1 (XNOR_4_1_NAND5_NUM725_OUT), .A2 (XNOR_4_2_NAND5_NUM725_OUT));

      NOR2_X1 XNOR_5_1_NAND5_NUM725 (.ZN (N2597), .A1 (XNOR_4_3_NAND5_NUM725_OUT), .A2 (GND));
      wire XNOR_1_1_NAND5_NUM726_OUT, XNOR_1_2_NAND5_NUM726_OUT, XNOR_1_3_NAND5_NUM726_OUT;
      NOR2_X1 XNOR_1_1_NAND5_NUM726 (.ZN (XNOR_1_1_NAND5_NUM726_OUT), .A1 (N2297), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND5_NUM726 (.ZN (XNOR_1_2_NAND5_NUM726_OUT), .A1 (GND), .A2 (N2427));
      NOR2_X1 XNOR_1_3_NAND5_NUM726 (.ZN (XNOR_1_3_NAND5_NUM726_OUT), .A1 (XNOR_1_1_NAND5_NUM726_OUT), .A2 (XNOR_1_2_NAND5_NUM726_OUT));

      wire XNOR_2_1_NAND5_NUM726_OUT, XNOR_2_2_NAND5_NUM726_OUT, XNOR_2_3_NAND5_NUM726_OUT;
      NOR2_X1 XNOR_2_1_NAND5_NUM726 (.ZN (XNOR_2_1_NAND5_NUM726_OUT), .A1 (N2375), .A2 (GND));
      NOR2_X1 XNOR_2_2_NAND5_NUM726 (.ZN (XNOR_2_2_NAND5_NUM726_OUT), .A1 (GND), .A2 (N2104));
      NOR2_X1 XNOR_2_3_NAND5_NUM726 (.ZN (XNOR_2_3_NAND5_NUM726_OUT), .A1 (XNOR_2_1_NAND5_NUM726_OUT), .A2 (XNOR_2_2_NAND5_NUM726_OUT));

      wire XNOR_3_1_NAND5_NUM726_OUT, XNOR_3_2_NAND5_NUM726_OUT, XNOR_3_3_NAND5_NUM726_OUT;
      NOR2_X1 XNOR_3_1_NAND5_NUM726 (.ZN (XNOR_3_1_NAND5_NUM726_OUT), .A1 (XNOR_1_3_NAND5_NUM726_OUT), .A2 (GND));
      NOR2_X1 XNOR_3_2_NAND5_NUM726 (.ZN (XNOR_3_2_NAND5_NUM726_OUT), .A1 (GND), .A2 (XNOR_2_3_NAND5_NUM726_OUT));
      NOR2_X1 XNOR_3_3_NAND5_NUM726 (.ZN (XNOR_3_3_NAND5_NUM726_OUT), .A1 (XNOR_3_1_NAND5_NUM726_OUT), .A2 (XNOR_3_2_NAND5_NUM726_OUT));

      wire XNOR_4_1_NAND5_NUM726_OUT, XNOR_4_2_NAND5_NUM726_OUT, XNOR_4_3_NAND5_NUM726_OUT;
      NOR2_X1 XNOR_4_1_NAND5_NUM726 (.ZN (XNOR_4_1_NAND5_NUM726_OUT), .A1 (N1171), .A2 (GND));
      NOR2_X1 XNOR_4_2_NAND5_NUM726 (.ZN (XNOR_4_2_NAND5_NUM726_OUT), .A1 (GND), .A2 (XNOR_3_3_NAND5_NUM726_OUT));
      NOR2_X1 XNOR_4_3_NAND5_NUM726 (.ZN (XNOR_4_3_NAND5_NUM726_OUT), .A1 (XNOR_4_1_NAND5_NUM726_OUT), .A2 (XNOR_4_2_NAND5_NUM726_OUT));

      NOR2_X1 XNOR_5_1_NAND5_NUM726 (.ZN (N2600), .A1 (XNOR_4_3_NAND5_NUM726_OUT), .A2 (GND));
      wire XNOR_1_1_NAND5_NUM727_OUT, XNOR_1_2_NAND5_NUM727_OUT, XNOR_1_3_NAND5_NUM727_OUT;
      NOR2_X1 XNOR_1_1_NAND5_NUM727 (.ZN (XNOR_1_1_NAND5_NUM727_OUT), .A1 (N2297), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND5_NUM727 (.ZN (XNOR_1_2_NAND5_NUM727_OUT), .A1 (GND), .A2 (N2427));
      NOR2_X1 XNOR_1_3_NAND5_NUM727 (.ZN (XNOR_1_3_NAND5_NUM727_OUT), .A1 (XNOR_1_1_NAND5_NUM727_OUT), .A2 (XNOR_1_2_NAND5_NUM727_OUT));

      wire XNOR_2_1_NAND5_NUM727_OUT, XNOR_2_2_NAND5_NUM727_OUT, XNOR_2_3_NAND5_NUM727_OUT;
      NOR2_X1 XNOR_2_1_NAND5_NUM727 (.ZN (XNOR_2_1_NAND5_NUM727_OUT), .A1 (N2340), .A2 (GND));
      NOR2_X1 XNOR_2_2_NAND5_NUM727 (.ZN (XNOR_2_2_NAND5_NUM727_OUT), .A1 (GND), .A2 (N2143));
      NOR2_X1 XNOR_2_3_NAND5_NUM727 (.ZN (XNOR_2_3_NAND5_NUM727_OUT), .A1 (XNOR_2_1_NAND5_NUM727_OUT), .A2 (XNOR_2_2_NAND5_NUM727_OUT));

      wire XNOR_3_1_NAND5_NUM727_OUT, XNOR_3_2_NAND5_NUM727_OUT, XNOR_3_3_NAND5_NUM727_OUT;
      NOR2_X1 XNOR_3_1_NAND5_NUM727 (.ZN (XNOR_3_1_NAND5_NUM727_OUT), .A1 (XNOR_1_3_NAND5_NUM727_OUT), .A2 (GND));
      NOR2_X1 XNOR_3_2_NAND5_NUM727 (.ZN (XNOR_3_2_NAND5_NUM727_OUT), .A1 (GND), .A2 (XNOR_2_3_NAND5_NUM727_OUT));
      NOR2_X1 XNOR_3_3_NAND5_NUM727 (.ZN (XNOR_3_3_NAND5_NUM727_OUT), .A1 (XNOR_3_1_NAND5_NUM727_OUT), .A2 (XNOR_3_2_NAND5_NUM727_OUT));

      wire XNOR_4_1_NAND5_NUM727_OUT, XNOR_4_2_NAND5_NUM727_OUT, XNOR_4_3_NAND5_NUM727_OUT;
      NOR2_X1 XNOR_4_1_NAND5_NUM727 (.ZN (XNOR_4_1_NAND5_NUM727_OUT), .A1 (N1171), .A2 (GND));
      NOR2_X1 XNOR_4_2_NAND5_NUM727 (.ZN (XNOR_4_2_NAND5_NUM727_OUT), .A1 (GND), .A2 (XNOR_3_3_NAND5_NUM727_OUT));
      NOR2_X1 XNOR_4_3_NAND5_NUM727 (.ZN (XNOR_4_3_NAND5_NUM727_OUT), .A1 (XNOR_4_1_NAND5_NUM727_OUT), .A2 (XNOR_4_2_NAND5_NUM727_OUT));

      NOR2_X1 XNOR_5_1_NAND5_NUM727 (.ZN (N2603), .A1 (XNOR_4_3_NAND5_NUM727_OUT), .A2 (GND));
      wire XNOR_1_1_NAND5_NUM728_OUT, XNOR_1_2_NAND5_NUM728_OUT, XNOR_1_3_NAND5_NUM728_OUT;
      NOR2_X1 XNOR_1_1_NAND5_NUM728 (.ZN (XNOR_1_1_NAND5_NUM728_OUT), .A1 (N2297), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND5_NUM728 (.ZN (XNOR_1_2_NAND5_NUM728_OUT), .A1 (GND), .A2 (N2427));
      NOR2_X1 XNOR_1_3_NAND5_NUM728 (.ZN (XNOR_1_3_NAND5_NUM728_OUT), .A1 (XNOR_1_1_NAND5_NUM728_OUT), .A2 (XNOR_1_2_NAND5_NUM728_OUT));

      wire XNOR_2_1_NAND5_NUM728_OUT, XNOR_2_2_NAND5_NUM728_OUT, XNOR_2_3_NAND5_NUM728_OUT;
      NOR2_X1 XNOR_2_1_NAND5_NUM728 (.ZN (XNOR_2_1_NAND5_NUM728_OUT), .A1 (N2353), .A2 (GND));
      NOR2_X1 XNOR_2_2_NAND5_NUM728 (.ZN (XNOR_2_2_NAND5_NUM728_OUT), .A1 (GND), .A2 (N2129));
      NOR2_X1 XNOR_2_3_NAND5_NUM728 (.ZN (XNOR_2_3_NAND5_NUM728_OUT), .A1 (XNOR_2_1_NAND5_NUM728_OUT), .A2 (XNOR_2_2_NAND5_NUM728_OUT));

      wire XNOR_3_1_NAND5_NUM728_OUT, XNOR_3_2_NAND5_NUM728_OUT, XNOR_3_3_NAND5_NUM728_OUT;
      NOR2_X1 XNOR_3_1_NAND5_NUM728 (.ZN (XNOR_3_1_NAND5_NUM728_OUT), .A1 (XNOR_1_3_NAND5_NUM728_OUT), .A2 (GND));
      NOR2_X1 XNOR_3_2_NAND5_NUM728 (.ZN (XNOR_3_2_NAND5_NUM728_OUT), .A1 (GND), .A2 (XNOR_2_3_NAND5_NUM728_OUT));
      NOR2_X1 XNOR_3_3_NAND5_NUM728 (.ZN (XNOR_3_3_NAND5_NUM728_OUT), .A1 (XNOR_3_1_NAND5_NUM728_OUT), .A2 (XNOR_3_2_NAND5_NUM728_OUT));

      wire XNOR_4_1_NAND5_NUM728_OUT, XNOR_4_2_NAND5_NUM728_OUT, XNOR_4_3_NAND5_NUM728_OUT;
      NOR2_X1 XNOR_4_1_NAND5_NUM728 (.ZN (XNOR_4_1_NAND5_NUM728_OUT), .A1 (N1188), .A2 (GND));
      NOR2_X1 XNOR_4_2_NAND5_NUM728 (.ZN (XNOR_4_2_NAND5_NUM728_OUT), .A1 (GND), .A2 (XNOR_3_3_NAND5_NUM728_OUT));
      NOR2_X1 XNOR_4_3_NAND5_NUM728 (.ZN (XNOR_4_3_NAND5_NUM728_OUT), .A1 (XNOR_4_1_NAND5_NUM728_OUT), .A2 (XNOR_4_2_NAND5_NUM728_OUT));

      NOR2_X1 XNOR_5_1_NAND5_NUM728 (.ZN (N2606), .A1 (XNOR_4_3_NAND5_NUM728_OUT), .A2 (GND));
      wire XNOR_1_1_NAND5_NUM729_OUT, XNOR_1_2_NAND5_NUM729_OUT, XNOR_1_3_NAND5_NUM729_OUT;
      NOR2_X1 XNOR_1_1_NAND5_NUM729 (.ZN (XNOR_1_1_NAND5_NUM729_OUT), .A1 (N2386), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND5_NUM729 (.ZN (XNOR_1_2_NAND5_NUM729_OUT), .A1 (GND), .A2 (N2326));
      NOR2_X1 XNOR_1_3_NAND5_NUM729 (.ZN (XNOR_1_3_NAND5_NUM729_OUT), .A1 (XNOR_1_1_NAND5_NUM729_OUT), .A2 (XNOR_1_2_NAND5_NUM729_OUT));

      wire XNOR_2_1_NAND5_NUM729_OUT, XNOR_2_2_NAND5_NUM729_OUT, XNOR_2_3_NAND5_NUM729_OUT;
      NOR2_X1 XNOR_2_1_NAND5_NUM729 (.ZN (XNOR_2_1_NAND5_NUM729_OUT), .A1 (N2361), .A2 (GND));
      NOR2_X1 XNOR_2_2_NAND5_NUM729 (.ZN (XNOR_2_2_NAND5_NUM729_OUT), .A1 (GND), .A2 (N2129));
      NOR2_X1 XNOR_2_3_NAND5_NUM729 (.ZN (XNOR_2_3_NAND5_NUM729_OUT), .A1 (XNOR_2_1_NAND5_NUM729_OUT), .A2 (XNOR_2_2_NAND5_NUM729_OUT));

      wire XNOR_3_1_NAND5_NUM729_OUT, XNOR_3_2_NAND5_NUM729_OUT, XNOR_3_3_NAND5_NUM729_OUT;
      NOR2_X1 XNOR_3_1_NAND5_NUM729 (.ZN (XNOR_3_1_NAND5_NUM729_OUT), .A1 (XNOR_1_3_NAND5_NUM729_OUT), .A2 (GND));
      NOR2_X1 XNOR_3_2_NAND5_NUM729 (.ZN (XNOR_3_2_NAND5_NUM729_OUT), .A1 (GND), .A2 (XNOR_2_3_NAND5_NUM729_OUT));
      NOR2_X1 XNOR_3_3_NAND5_NUM729 (.ZN (XNOR_3_3_NAND5_NUM729_OUT), .A1 (XNOR_3_1_NAND5_NUM729_OUT), .A2 (XNOR_3_2_NAND5_NUM729_OUT));

      wire XNOR_4_1_NAND5_NUM729_OUT, XNOR_4_2_NAND5_NUM729_OUT, XNOR_4_3_NAND5_NUM729_OUT;
      NOR2_X1 XNOR_4_1_NAND5_NUM729 (.ZN (XNOR_4_1_NAND5_NUM729_OUT), .A1 (N1188), .A2 (GND));
      NOR2_X1 XNOR_4_2_NAND5_NUM729 (.ZN (XNOR_4_2_NAND5_NUM729_OUT), .A1 (GND), .A2 (XNOR_3_3_NAND5_NUM729_OUT));
      NOR2_X1 XNOR_4_3_NAND5_NUM729 (.ZN (XNOR_4_3_NAND5_NUM729_OUT), .A1 (XNOR_4_1_NAND5_NUM729_OUT), .A2 (XNOR_4_2_NAND5_NUM729_OUT));

      NOR2_X1 XNOR_5_1_NAND5_NUM729 (.ZN (N2611), .A1 (XNOR_4_3_NAND5_NUM729_OUT), .A2 (GND));
      wire XNOR_1_1_NAND5_NUM730_OUT, XNOR_1_2_NAND5_NUM730_OUT, XNOR_1_3_NAND5_NUM730_OUT;
      NOR2_X1 XNOR_1_1_NAND5_NUM730 (.ZN (XNOR_1_1_NAND5_NUM730_OUT), .A1 (N2386), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND5_NUM730 (.ZN (XNOR_1_2_NAND5_NUM730_OUT), .A1 (GND), .A2 (N2326));
      NOR2_X1 XNOR_1_3_NAND5_NUM730 (.ZN (XNOR_1_3_NAND5_NUM730_OUT), .A1 (XNOR_1_1_NAND5_NUM730_OUT), .A2 (XNOR_1_2_NAND5_NUM730_OUT));

      wire XNOR_2_1_NAND5_NUM730_OUT, XNOR_2_2_NAND5_NUM730_OUT, XNOR_2_3_NAND5_NUM730_OUT;
      NOR2_X1 XNOR_2_1_NAND5_NUM730 (.ZN (XNOR_2_1_NAND5_NUM730_OUT), .A1 (N2361), .A2 (GND));
      NOR2_X1 XNOR_2_2_NAND5_NUM730 (.ZN (XNOR_2_2_NAND5_NUM730_OUT), .A1 (GND), .A2 (N2119));
      NOR2_X1 XNOR_2_3_NAND5_NUM730 (.ZN (XNOR_2_3_NAND5_NUM730_OUT), .A1 (XNOR_2_1_NAND5_NUM730_OUT), .A2 (XNOR_2_2_NAND5_NUM730_OUT));

      wire XNOR_3_1_NAND5_NUM730_OUT, XNOR_3_2_NAND5_NUM730_OUT, XNOR_3_3_NAND5_NUM730_OUT;
      NOR2_X1 XNOR_3_1_NAND5_NUM730 (.ZN (XNOR_3_1_NAND5_NUM730_OUT), .A1 (XNOR_1_3_NAND5_NUM730_OUT), .A2 (GND));
      NOR2_X1 XNOR_3_2_NAND5_NUM730 (.ZN (XNOR_3_2_NAND5_NUM730_OUT), .A1 (GND), .A2 (XNOR_2_3_NAND5_NUM730_OUT));
      NOR2_X1 XNOR_3_3_NAND5_NUM730 (.ZN (XNOR_3_3_NAND5_NUM730_OUT), .A1 (XNOR_3_1_NAND5_NUM730_OUT), .A2 (XNOR_3_2_NAND5_NUM730_OUT));

      wire XNOR_4_1_NAND5_NUM730_OUT, XNOR_4_2_NAND5_NUM730_OUT, XNOR_4_3_NAND5_NUM730_OUT;
      NOR2_X1 XNOR_4_1_NAND5_NUM730 (.ZN (XNOR_4_1_NAND5_NUM730_OUT), .A1 (N1188), .A2 (GND));
      NOR2_X1 XNOR_4_2_NAND5_NUM730 (.ZN (XNOR_4_2_NAND5_NUM730_OUT), .A1 (GND), .A2 (XNOR_3_3_NAND5_NUM730_OUT));
      NOR2_X1 XNOR_4_3_NAND5_NUM730 (.ZN (XNOR_4_3_NAND5_NUM730_OUT), .A1 (XNOR_4_1_NAND5_NUM730_OUT), .A2 (XNOR_4_2_NAND5_NUM730_OUT));

      NOR2_X1 XNOR_5_1_NAND5_NUM730 (.ZN (N2614), .A1 (XNOR_4_3_NAND5_NUM730_OUT), .A2 (GND));
      wire XNOR_1_1_NAND5_NUM731_OUT, XNOR_1_2_NAND5_NUM731_OUT, XNOR_1_3_NAND5_NUM731_OUT;
      NOR2_X1 XNOR_1_1_NAND5_NUM731 (.ZN (XNOR_1_1_NAND5_NUM731_OUT), .A1 (N2386), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND5_NUM731 (.ZN (XNOR_1_2_NAND5_NUM731_OUT), .A1 (GND), .A2 (N2326));
      NOR2_X1 XNOR_1_3_NAND5_NUM731 (.ZN (XNOR_1_3_NAND5_NUM731_OUT), .A1 (XNOR_1_1_NAND5_NUM731_OUT), .A2 (XNOR_1_2_NAND5_NUM731_OUT));

      wire XNOR_2_1_NAND5_NUM731_OUT, XNOR_2_2_NAND5_NUM731_OUT, XNOR_2_3_NAND5_NUM731_OUT;
      NOR2_X1 XNOR_2_1_NAND5_NUM731 (.ZN (XNOR_2_1_NAND5_NUM731_OUT), .A1 (N2375), .A2 (GND));
      NOR2_X1 XNOR_2_2_NAND5_NUM731 (.ZN (XNOR_2_2_NAND5_NUM731_OUT), .A1 (GND), .A2 (N2104));
      NOR2_X1 XNOR_2_3_NAND5_NUM731 (.ZN (XNOR_2_3_NAND5_NUM731_OUT), .A1 (XNOR_2_1_NAND5_NUM731_OUT), .A2 (XNOR_2_2_NAND5_NUM731_OUT));

      wire XNOR_3_1_NAND5_NUM731_OUT, XNOR_3_2_NAND5_NUM731_OUT, XNOR_3_3_NAND5_NUM731_OUT;
      NOR2_X1 XNOR_3_1_NAND5_NUM731 (.ZN (XNOR_3_1_NAND5_NUM731_OUT), .A1 (XNOR_1_3_NAND5_NUM731_OUT), .A2 (GND));
      NOR2_X1 XNOR_3_2_NAND5_NUM731 (.ZN (XNOR_3_2_NAND5_NUM731_OUT), .A1 (GND), .A2 (XNOR_2_3_NAND5_NUM731_OUT));
      NOR2_X1 XNOR_3_3_NAND5_NUM731 (.ZN (XNOR_3_3_NAND5_NUM731_OUT), .A1 (XNOR_3_1_NAND5_NUM731_OUT), .A2 (XNOR_3_2_NAND5_NUM731_OUT));

      wire XNOR_4_1_NAND5_NUM731_OUT, XNOR_4_2_NAND5_NUM731_OUT, XNOR_4_3_NAND5_NUM731_OUT;
      NOR2_X1 XNOR_4_1_NAND5_NUM731 (.ZN (XNOR_4_1_NAND5_NUM731_OUT), .A1 (N1188), .A2 (GND));
      NOR2_X1 XNOR_4_2_NAND5_NUM731 (.ZN (XNOR_4_2_NAND5_NUM731_OUT), .A1 (GND), .A2 (XNOR_3_3_NAND5_NUM731_OUT));
      NOR2_X1 XNOR_4_3_NAND5_NUM731 (.ZN (XNOR_4_3_NAND5_NUM731_OUT), .A1 (XNOR_4_1_NAND5_NUM731_OUT), .A2 (XNOR_4_2_NAND5_NUM731_OUT));

      NOR2_X1 XNOR_5_1_NAND5_NUM731 (.ZN (N2617), .A1 (XNOR_4_3_NAND5_NUM731_OUT), .A2 (GND));
      wire XNOR_1_1_NAND5_NUM732_OUT, XNOR_1_2_NAND5_NUM732_OUT, XNOR_1_3_NAND5_NUM732_OUT;
      NOR2_X1 XNOR_1_1_NAND5_NUM732 (.ZN (XNOR_1_1_NAND5_NUM732_OUT), .A1 (N2386), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND5_NUM732 (.ZN (XNOR_1_2_NAND5_NUM732_OUT), .A1 (GND), .A2 (N2326));
      NOR2_X1 XNOR_1_3_NAND5_NUM732 (.ZN (XNOR_1_3_NAND5_NUM732_OUT), .A1 (XNOR_1_1_NAND5_NUM732_OUT), .A2 (XNOR_1_2_NAND5_NUM732_OUT));

      wire XNOR_2_1_NAND5_NUM732_OUT, XNOR_2_2_NAND5_NUM732_OUT, XNOR_2_3_NAND5_NUM732_OUT;
      NOR2_X1 XNOR_2_1_NAND5_NUM732 (.ZN (XNOR_2_1_NAND5_NUM732_OUT), .A1 (N2353), .A2 (GND));
      NOR2_X1 XNOR_2_2_NAND5_NUM732 (.ZN (XNOR_2_2_NAND5_NUM732_OUT), .A1 (GND), .A2 (N2129));
      NOR2_X1 XNOR_2_3_NAND5_NUM732 (.ZN (XNOR_2_3_NAND5_NUM732_OUT), .A1 (XNOR_2_1_NAND5_NUM732_OUT), .A2 (XNOR_2_2_NAND5_NUM732_OUT));

      wire XNOR_3_1_NAND5_NUM732_OUT, XNOR_3_2_NAND5_NUM732_OUT, XNOR_3_3_NAND5_NUM732_OUT;
      NOR2_X1 XNOR_3_1_NAND5_NUM732 (.ZN (XNOR_3_1_NAND5_NUM732_OUT), .A1 (XNOR_1_3_NAND5_NUM732_OUT), .A2 (GND));
      NOR2_X1 XNOR_3_2_NAND5_NUM732 (.ZN (XNOR_3_2_NAND5_NUM732_OUT), .A1 (GND), .A2 (XNOR_2_3_NAND5_NUM732_OUT));
      NOR2_X1 XNOR_3_3_NAND5_NUM732 (.ZN (XNOR_3_3_NAND5_NUM732_OUT), .A1 (XNOR_3_1_NAND5_NUM732_OUT), .A2 (XNOR_3_2_NAND5_NUM732_OUT));

      wire XNOR_4_1_NAND5_NUM732_OUT, XNOR_4_2_NAND5_NUM732_OUT, XNOR_4_3_NAND5_NUM732_OUT;
      NOR2_X1 XNOR_4_1_NAND5_NUM732 (.ZN (XNOR_4_1_NAND5_NUM732_OUT), .A1 (N1188), .A2 (GND));
      NOR2_X1 XNOR_4_2_NAND5_NUM732 (.ZN (XNOR_4_2_NAND5_NUM732_OUT), .A1 (GND), .A2 (XNOR_3_3_NAND5_NUM732_OUT));
      NOR2_X1 XNOR_4_3_NAND5_NUM732 (.ZN (XNOR_4_3_NAND5_NUM732_OUT), .A1 (XNOR_4_1_NAND5_NUM732_OUT), .A2 (XNOR_4_2_NAND5_NUM732_OUT));

      NOR2_X1 XNOR_5_1_NAND5_NUM732 (.ZN (N2620), .A1 (XNOR_4_3_NAND5_NUM732_OUT), .A2 (GND));
      wire XNOR_1_1_NAND5_NUM733_OUT, XNOR_1_2_NAND5_NUM733_OUT, XNOR_1_3_NAND5_NUM733_OUT;
      NOR2_X1 XNOR_1_1_NAND5_NUM733 (.ZN (XNOR_1_1_NAND5_NUM733_OUT), .A1 (N2297), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND5_NUM733 (.ZN (XNOR_1_2_NAND5_NUM733_OUT), .A1 (GND), .A2 (N2427));
      NOR2_X1 XNOR_1_3_NAND5_NUM733 (.ZN (XNOR_1_3_NAND5_NUM733_OUT), .A1 (XNOR_1_1_NAND5_NUM733_OUT), .A2 (XNOR_1_2_NAND5_NUM733_OUT));

      wire XNOR_2_1_NAND5_NUM733_OUT, XNOR_2_2_NAND5_NUM733_OUT, XNOR_2_3_NAND5_NUM733_OUT;
      NOR2_X1 XNOR_2_1_NAND5_NUM733 (.ZN (XNOR_2_1_NAND5_NUM733_OUT), .A1 (N2340), .A2 (GND));
      NOR2_X1 XNOR_2_2_NAND5_NUM733 (.ZN (XNOR_2_2_NAND5_NUM733_OUT), .A1 (GND), .A2 (N2104));
      NOR2_X1 XNOR_2_3_NAND5_NUM733 (.ZN (XNOR_2_3_NAND5_NUM733_OUT), .A1 (XNOR_2_1_NAND5_NUM733_OUT), .A2 (XNOR_2_2_NAND5_NUM733_OUT));

      wire XNOR_3_1_NAND5_NUM733_OUT, XNOR_3_2_NAND5_NUM733_OUT, XNOR_3_3_NAND5_NUM733_OUT;
      NOR2_X1 XNOR_3_1_NAND5_NUM733 (.ZN (XNOR_3_1_NAND5_NUM733_OUT), .A1 (XNOR_1_3_NAND5_NUM733_OUT), .A2 (GND));
      NOR2_X1 XNOR_3_2_NAND5_NUM733 (.ZN (XNOR_3_2_NAND5_NUM733_OUT), .A1 (GND), .A2 (XNOR_2_3_NAND5_NUM733_OUT));
      NOR2_X1 XNOR_3_3_NAND5_NUM733 (.ZN (XNOR_3_3_NAND5_NUM733_OUT), .A1 (XNOR_3_1_NAND5_NUM733_OUT), .A2 (XNOR_3_2_NAND5_NUM733_OUT));

      wire XNOR_4_1_NAND5_NUM733_OUT, XNOR_4_2_NAND5_NUM733_OUT, XNOR_4_3_NAND5_NUM733_OUT;
      NOR2_X1 XNOR_4_1_NAND5_NUM733 (.ZN (XNOR_4_1_NAND5_NUM733_OUT), .A1 (N926), .A2 (GND));
      NOR2_X1 XNOR_4_2_NAND5_NUM733 (.ZN (XNOR_4_2_NAND5_NUM733_OUT), .A1 (GND), .A2 (XNOR_3_3_NAND5_NUM733_OUT));
      NOR2_X1 XNOR_4_3_NAND5_NUM733 (.ZN (XNOR_4_3_NAND5_NUM733_OUT), .A1 (XNOR_4_1_NAND5_NUM733_OUT), .A2 (XNOR_4_2_NAND5_NUM733_OUT));

      NOR2_X1 XNOR_5_1_NAND5_NUM733 (.ZN (N2627), .A1 (XNOR_4_3_NAND5_NUM733_OUT), .A2 (GND));
      wire XNOR_1_1_NAND5_NUM734_OUT, XNOR_1_2_NAND5_NUM734_OUT, XNOR_1_3_NAND5_NUM734_OUT;
      NOR2_X1 XNOR_1_1_NAND5_NUM734 (.ZN (XNOR_1_1_NAND5_NUM734_OUT), .A1 (N2386), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND5_NUM734 (.ZN (XNOR_1_2_NAND5_NUM734_OUT), .A1 (GND), .A2 (N2326));
      NOR2_X1 XNOR_1_3_NAND5_NUM734 (.ZN (XNOR_1_3_NAND5_NUM734_OUT), .A1 (XNOR_1_1_NAND5_NUM734_OUT), .A2 (XNOR_1_2_NAND5_NUM734_OUT));

      wire XNOR_2_1_NAND5_NUM734_OUT, XNOR_2_2_NAND5_NUM734_OUT, XNOR_2_3_NAND5_NUM734_OUT;
      NOR2_X1 XNOR_2_1_NAND5_NUM734 (.ZN (XNOR_2_1_NAND5_NUM734_OUT), .A1 (N2340), .A2 (GND));
      NOR2_X1 XNOR_2_2_NAND5_NUM734 (.ZN (XNOR_2_2_NAND5_NUM734_OUT), .A1 (GND), .A2 (N2104));
      NOR2_X1 XNOR_2_3_NAND5_NUM734 (.ZN (XNOR_2_3_NAND5_NUM734_OUT), .A1 (XNOR_2_1_NAND5_NUM734_OUT), .A2 (XNOR_2_2_NAND5_NUM734_OUT));

      wire XNOR_3_1_NAND5_NUM734_OUT, XNOR_3_2_NAND5_NUM734_OUT, XNOR_3_3_NAND5_NUM734_OUT;
      NOR2_X1 XNOR_3_1_NAND5_NUM734 (.ZN (XNOR_3_1_NAND5_NUM734_OUT), .A1 (XNOR_1_3_NAND5_NUM734_OUT), .A2 (GND));
      NOR2_X1 XNOR_3_2_NAND5_NUM734 (.ZN (XNOR_3_2_NAND5_NUM734_OUT), .A1 (GND), .A2 (XNOR_2_3_NAND5_NUM734_OUT));
      NOR2_X1 XNOR_3_3_NAND5_NUM734 (.ZN (XNOR_3_3_NAND5_NUM734_OUT), .A1 (XNOR_3_1_NAND5_NUM734_OUT), .A2 (XNOR_3_2_NAND5_NUM734_OUT));

      wire XNOR_4_1_NAND5_NUM734_OUT, XNOR_4_2_NAND5_NUM734_OUT, XNOR_4_3_NAND5_NUM734_OUT;
      NOR2_X1 XNOR_4_1_NAND5_NUM734 (.ZN (XNOR_4_1_NAND5_NUM734_OUT), .A1 (N926), .A2 (GND));
      NOR2_X1 XNOR_4_2_NAND5_NUM734 (.ZN (XNOR_4_2_NAND5_NUM734_OUT), .A1 (GND), .A2 (XNOR_3_3_NAND5_NUM734_OUT));
      NOR2_X1 XNOR_4_3_NAND5_NUM734 (.ZN (XNOR_4_3_NAND5_NUM734_OUT), .A1 (XNOR_4_1_NAND5_NUM734_OUT), .A2 (XNOR_4_2_NAND5_NUM734_OUT));

      NOR2_X1 XNOR_5_1_NAND5_NUM734 (.ZN (N2628), .A1 (XNOR_4_3_NAND5_NUM734_OUT), .A2 (GND));
      wire XNOR_1_1_NAND5_NUM735_OUT, XNOR_1_2_NAND5_NUM735_OUT, XNOR_1_3_NAND5_NUM735_OUT;
      NOR2_X1 XNOR_1_1_NAND5_NUM735 (.ZN (XNOR_1_1_NAND5_NUM735_OUT), .A1 (N2386), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND5_NUM735 (.ZN (XNOR_1_2_NAND5_NUM735_OUT), .A1 (GND), .A2 (N2427));
      NOR2_X1 XNOR_1_3_NAND5_NUM735 (.ZN (XNOR_1_3_NAND5_NUM735_OUT), .A1 (XNOR_1_1_NAND5_NUM735_OUT), .A2 (XNOR_1_2_NAND5_NUM735_OUT));

      wire XNOR_2_1_NAND5_NUM735_OUT, XNOR_2_2_NAND5_NUM735_OUT, XNOR_2_3_NAND5_NUM735_OUT;
      NOR2_X1 XNOR_2_1_NAND5_NUM735 (.ZN (XNOR_2_1_NAND5_NUM735_OUT), .A1 (N2361), .A2 (GND));
      NOR2_X1 XNOR_2_2_NAND5_NUM735 (.ZN (XNOR_2_2_NAND5_NUM735_OUT), .A1 (GND), .A2 (N2104));
      NOR2_X1 XNOR_2_3_NAND5_NUM735 (.ZN (XNOR_2_3_NAND5_NUM735_OUT), .A1 (XNOR_2_1_NAND5_NUM735_OUT), .A2 (XNOR_2_2_NAND5_NUM735_OUT));

      wire XNOR_3_1_NAND5_NUM735_OUT, XNOR_3_2_NAND5_NUM735_OUT, XNOR_3_3_NAND5_NUM735_OUT;
      NOR2_X1 XNOR_3_1_NAND5_NUM735 (.ZN (XNOR_3_1_NAND5_NUM735_OUT), .A1 (XNOR_1_3_NAND5_NUM735_OUT), .A2 (GND));
      NOR2_X1 XNOR_3_2_NAND5_NUM735 (.ZN (XNOR_3_2_NAND5_NUM735_OUT), .A1 (GND), .A2 (XNOR_2_3_NAND5_NUM735_OUT));
      NOR2_X1 XNOR_3_3_NAND5_NUM735 (.ZN (XNOR_3_3_NAND5_NUM735_OUT), .A1 (XNOR_3_1_NAND5_NUM735_OUT), .A2 (XNOR_3_2_NAND5_NUM735_OUT));

      wire XNOR_4_1_NAND5_NUM735_OUT, XNOR_4_2_NAND5_NUM735_OUT, XNOR_4_3_NAND5_NUM735_OUT;
      NOR2_X1 XNOR_4_1_NAND5_NUM735 (.ZN (XNOR_4_1_NAND5_NUM735_OUT), .A1 (N926), .A2 (GND));
      NOR2_X1 XNOR_4_2_NAND5_NUM735 (.ZN (XNOR_4_2_NAND5_NUM735_OUT), .A1 (GND), .A2 (XNOR_3_3_NAND5_NUM735_OUT));
      NOR2_X1 XNOR_4_3_NAND5_NUM735 (.ZN (XNOR_4_3_NAND5_NUM735_OUT), .A1 (XNOR_4_1_NAND5_NUM735_OUT), .A2 (XNOR_4_2_NAND5_NUM735_OUT));

      NOR2_X1 XNOR_5_1_NAND5_NUM735 (.ZN (N2629), .A1 (XNOR_4_3_NAND5_NUM735_OUT), .A2 (GND));
      wire XNOR_1_1_NAND5_NUM736_OUT, XNOR_1_2_NAND5_NUM736_OUT, XNOR_1_3_NAND5_NUM736_OUT;
      NOR2_X1 XNOR_1_1_NAND5_NUM736 (.ZN (XNOR_1_1_NAND5_NUM736_OUT), .A1 (N2386), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND5_NUM736 (.ZN (XNOR_1_2_NAND5_NUM736_OUT), .A1 (GND), .A2 (N2427));
      NOR2_X1 XNOR_1_3_NAND5_NUM736 (.ZN (XNOR_1_3_NAND5_NUM736_OUT), .A1 (XNOR_1_1_NAND5_NUM736_OUT), .A2 (XNOR_1_2_NAND5_NUM736_OUT));

      wire XNOR_2_1_NAND5_NUM736_OUT, XNOR_2_2_NAND5_NUM736_OUT, XNOR_2_3_NAND5_NUM736_OUT;
      NOR2_X1 XNOR_2_1_NAND5_NUM736 (.ZN (XNOR_2_1_NAND5_NUM736_OUT), .A1 (N2340), .A2 (GND));
      NOR2_X1 XNOR_2_2_NAND5_NUM736 (.ZN (XNOR_2_2_NAND5_NUM736_OUT), .A1 (GND), .A2 (N2129));
      NOR2_X1 XNOR_2_3_NAND5_NUM736 (.ZN (XNOR_2_3_NAND5_NUM736_OUT), .A1 (XNOR_2_1_NAND5_NUM736_OUT), .A2 (XNOR_2_2_NAND5_NUM736_OUT));

      wire XNOR_3_1_NAND5_NUM736_OUT, XNOR_3_2_NAND5_NUM736_OUT, XNOR_3_3_NAND5_NUM736_OUT;
      NOR2_X1 XNOR_3_1_NAND5_NUM736 (.ZN (XNOR_3_1_NAND5_NUM736_OUT), .A1 (XNOR_1_3_NAND5_NUM736_OUT), .A2 (GND));
      NOR2_X1 XNOR_3_2_NAND5_NUM736 (.ZN (XNOR_3_2_NAND5_NUM736_OUT), .A1 (GND), .A2 (XNOR_2_3_NAND5_NUM736_OUT));
      NOR2_X1 XNOR_3_3_NAND5_NUM736 (.ZN (XNOR_3_3_NAND5_NUM736_OUT), .A1 (XNOR_3_1_NAND5_NUM736_OUT), .A2 (XNOR_3_2_NAND5_NUM736_OUT));

      wire XNOR_4_1_NAND5_NUM736_OUT, XNOR_4_2_NAND5_NUM736_OUT, XNOR_4_3_NAND5_NUM736_OUT;
      NOR2_X1 XNOR_4_1_NAND5_NUM736 (.ZN (XNOR_4_1_NAND5_NUM736_OUT), .A1 (N926), .A2 (GND));
      NOR2_X1 XNOR_4_2_NAND5_NUM736 (.ZN (XNOR_4_2_NAND5_NUM736_OUT), .A1 (GND), .A2 (XNOR_3_3_NAND5_NUM736_OUT));
      NOR2_X1 XNOR_4_3_NAND5_NUM736 (.ZN (XNOR_4_3_NAND5_NUM736_OUT), .A1 (XNOR_4_1_NAND5_NUM736_OUT), .A2 (XNOR_4_2_NAND5_NUM736_OUT));

      NOR2_X1 XNOR_5_1_NAND5_NUM736 (.ZN (N2630), .A1 (XNOR_4_3_NAND5_NUM736_OUT), .A2 (GND));
      wire XNOR_1_1_NAND5_NUM737_OUT, XNOR_1_2_NAND5_NUM737_OUT, XNOR_1_3_NAND5_NUM737_OUT;
      NOR2_X1 XNOR_1_1_NAND5_NUM737 (.ZN (XNOR_1_1_NAND5_NUM737_OUT), .A1 (N2386), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND5_NUM737 (.ZN (XNOR_1_2_NAND5_NUM737_OUT), .A1 (GND), .A2 (N2427));
      NOR2_X1 XNOR_1_3_NAND5_NUM737 (.ZN (XNOR_1_3_NAND5_NUM737_OUT), .A1 (XNOR_1_1_NAND5_NUM737_OUT), .A2 (XNOR_1_2_NAND5_NUM737_OUT));

      wire XNOR_2_1_NAND5_NUM737_OUT, XNOR_2_2_NAND5_NUM737_OUT, XNOR_2_3_NAND5_NUM737_OUT;
      NOR2_X1 XNOR_2_1_NAND5_NUM737 (.ZN (XNOR_2_1_NAND5_NUM737_OUT), .A1 (N2340), .A2 (GND));
      NOR2_X1 XNOR_2_2_NAND5_NUM737 (.ZN (XNOR_2_2_NAND5_NUM737_OUT), .A1 (GND), .A2 (N2119));
      NOR2_X1 XNOR_2_3_NAND5_NUM737 (.ZN (XNOR_2_3_NAND5_NUM737_OUT), .A1 (XNOR_2_1_NAND5_NUM737_OUT), .A2 (XNOR_2_2_NAND5_NUM737_OUT));

      wire XNOR_3_1_NAND5_NUM737_OUT, XNOR_3_2_NAND5_NUM737_OUT, XNOR_3_3_NAND5_NUM737_OUT;
      NOR2_X1 XNOR_3_1_NAND5_NUM737 (.ZN (XNOR_3_1_NAND5_NUM737_OUT), .A1 (XNOR_1_3_NAND5_NUM737_OUT), .A2 (GND));
      NOR2_X1 XNOR_3_2_NAND5_NUM737 (.ZN (XNOR_3_2_NAND5_NUM737_OUT), .A1 (GND), .A2 (XNOR_2_3_NAND5_NUM737_OUT));
      NOR2_X1 XNOR_3_3_NAND5_NUM737 (.ZN (XNOR_3_3_NAND5_NUM737_OUT), .A1 (XNOR_3_1_NAND5_NUM737_OUT), .A2 (XNOR_3_2_NAND5_NUM737_OUT));

      wire XNOR_4_1_NAND5_NUM737_OUT, XNOR_4_2_NAND5_NUM737_OUT, XNOR_4_3_NAND5_NUM737_OUT;
      NOR2_X1 XNOR_4_1_NAND5_NUM737 (.ZN (XNOR_4_1_NAND5_NUM737_OUT), .A1 (N926), .A2 (GND));
      NOR2_X1 XNOR_4_2_NAND5_NUM737 (.ZN (XNOR_4_2_NAND5_NUM737_OUT), .A1 (GND), .A2 (XNOR_3_3_NAND5_NUM737_OUT));
      NOR2_X1 XNOR_4_3_NAND5_NUM737 (.ZN (XNOR_4_3_NAND5_NUM737_OUT), .A1 (XNOR_4_1_NAND5_NUM737_OUT), .A2 (XNOR_4_2_NAND5_NUM737_OUT));

      NOR2_X1 XNOR_5_1_NAND5_NUM737 (.ZN (N2631), .A1 (XNOR_4_3_NAND5_NUM737_OUT), .A2 (GND));
      wire XNOR_1_1_NAND5_NUM738_OUT, XNOR_1_2_NAND5_NUM738_OUT, XNOR_1_3_NAND5_NUM738_OUT;
      NOR2_X1 XNOR_1_1_NAND5_NUM738 (.ZN (XNOR_1_1_NAND5_NUM738_OUT), .A1 (N2386), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND5_NUM738 (.ZN (XNOR_1_2_NAND5_NUM738_OUT), .A1 (GND), .A2 (N2427));
      NOR2_X1 XNOR_1_3_NAND5_NUM738 (.ZN (XNOR_1_3_NAND5_NUM738_OUT), .A1 (XNOR_1_1_NAND5_NUM738_OUT), .A2 (XNOR_1_2_NAND5_NUM738_OUT));

      wire XNOR_2_1_NAND5_NUM738_OUT, XNOR_2_2_NAND5_NUM738_OUT, XNOR_2_3_NAND5_NUM738_OUT;
      NOR2_X1 XNOR_2_1_NAND5_NUM738 (.ZN (XNOR_2_1_NAND5_NUM738_OUT), .A1 (N2353), .A2 (GND));
      NOR2_X1 XNOR_2_2_NAND5_NUM738 (.ZN (XNOR_2_2_NAND5_NUM738_OUT), .A1 (GND), .A2 (N2104));
      NOR2_X1 XNOR_2_3_NAND5_NUM738 (.ZN (XNOR_2_3_NAND5_NUM738_OUT), .A1 (XNOR_2_1_NAND5_NUM738_OUT), .A2 (XNOR_2_2_NAND5_NUM738_OUT));

      wire XNOR_3_1_NAND5_NUM738_OUT, XNOR_3_2_NAND5_NUM738_OUT, XNOR_3_3_NAND5_NUM738_OUT;
      NOR2_X1 XNOR_3_1_NAND5_NUM738 (.ZN (XNOR_3_1_NAND5_NUM738_OUT), .A1 (XNOR_1_3_NAND5_NUM738_OUT), .A2 (GND));
      NOR2_X1 XNOR_3_2_NAND5_NUM738 (.ZN (XNOR_3_2_NAND5_NUM738_OUT), .A1 (GND), .A2 (XNOR_2_3_NAND5_NUM738_OUT));
      NOR2_X1 XNOR_3_3_NAND5_NUM738 (.ZN (XNOR_3_3_NAND5_NUM738_OUT), .A1 (XNOR_3_1_NAND5_NUM738_OUT), .A2 (XNOR_3_2_NAND5_NUM738_OUT));

      wire XNOR_4_1_NAND5_NUM738_OUT, XNOR_4_2_NAND5_NUM738_OUT, XNOR_4_3_NAND5_NUM738_OUT;
      NOR2_X1 XNOR_4_1_NAND5_NUM738 (.ZN (XNOR_4_1_NAND5_NUM738_OUT), .A1 (N926), .A2 (GND));
      NOR2_X1 XNOR_4_2_NAND5_NUM738 (.ZN (XNOR_4_2_NAND5_NUM738_OUT), .A1 (GND), .A2 (XNOR_3_3_NAND5_NUM738_OUT));
      NOR2_X1 XNOR_4_3_NAND5_NUM738 (.ZN (XNOR_4_3_NAND5_NUM738_OUT), .A1 (XNOR_4_1_NAND5_NUM738_OUT), .A2 (XNOR_4_2_NAND5_NUM738_OUT));

      NOR2_X1 XNOR_5_1_NAND5_NUM738 (.ZN (N2632), .A1 (XNOR_4_3_NAND5_NUM738_OUT), .A2 (GND));
      wire XNOR_1_1_NAND5_NUM739_OUT, XNOR_1_2_NAND5_NUM739_OUT, XNOR_1_3_NAND5_NUM739_OUT;
      NOR2_X1 XNOR_1_1_NAND5_NUM739 (.ZN (XNOR_1_1_NAND5_NUM739_OUT), .A1 (N2386), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND5_NUM739 (.ZN (XNOR_1_2_NAND5_NUM739_OUT), .A1 (GND), .A2 (N2426));
      NOR2_X1 XNOR_1_3_NAND5_NUM739 (.ZN (XNOR_1_3_NAND5_NUM739_OUT), .A1 (XNOR_1_1_NAND5_NUM739_OUT), .A2 (XNOR_1_2_NAND5_NUM739_OUT));

      wire XNOR_2_1_NAND5_NUM739_OUT, XNOR_2_2_NAND5_NUM739_OUT, XNOR_2_3_NAND5_NUM739_OUT;
      NOR2_X1 XNOR_2_1_NAND5_NUM739 (.ZN (XNOR_2_1_NAND5_NUM739_OUT), .A1 (N2340), .A2 (GND));
      NOR2_X1 XNOR_2_2_NAND5_NUM739 (.ZN (XNOR_2_2_NAND5_NUM739_OUT), .A1 (GND), .A2 (N2104));
      NOR2_X1 XNOR_2_3_NAND5_NUM739 (.ZN (XNOR_2_3_NAND5_NUM739_OUT), .A1 (XNOR_2_1_NAND5_NUM739_OUT), .A2 (XNOR_2_2_NAND5_NUM739_OUT));

      wire XNOR_3_1_NAND5_NUM739_OUT, XNOR_3_2_NAND5_NUM739_OUT, XNOR_3_3_NAND5_NUM739_OUT;
      NOR2_X1 XNOR_3_1_NAND5_NUM739 (.ZN (XNOR_3_1_NAND5_NUM739_OUT), .A1 (XNOR_1_3_NAND5_NUM739_OUT), .A2 (GND));
      NOR2_X1 XNOR_3_2_NAND5_NUM739 (.ZN (XNOR_3_2_NAND5_NUM739_OUT), .A1 (GND), .A2 (XNOR_2_3_NAND5_NUM739_OUT));
      NOR2_X1 XNOR_3_3_NAND5_NUM739 (.ZN (XNOR_3_3_NAND5_NUM739_OUT), .A1 (XNOR_3_1_NAND5_NUM739_OUT), .A2 (XNOR_3_2_NAND5_NUM739_OUT));

      wire XNOR_4_1_NAND5_NUM739_OUT, XNOR_4_2_NAND5_NUM739_OUT, XNOR_4_3_NAND5_NUM739_OUT;
      NOR2_X1 XNOR_4_1_NAND5_NUM739 (.ZN (XNOR_4_1_NAND5_NUM739_OUT), .A1 (N926), .A2 (GND));
      NOR2_X1 XNOR_4_2_NAND5_NUM739 (.ZN (XNOR_4_2_NAND5_NUM739_OUT), .A1 (GND), .A2 (XNOR_3_3_NAND5_NUM739_OUT));
      NOR2_X1 XNOR_4_3_NAND5_NUM739 (.ZN (XNOR_4_3_NAND5_NUM739_OUT), .A1 (XNOR_4_1_NAND5_NUM739_OUT), .A2 (XNOR_4_2_NAND5_NUM739_OUT));

      NOR2_X1 XNOR_5_1_NAND5_NUM739 (.ZN (N2633), .A1 (XNOR_4_3_NAND5_NUM739_OUT), .A2 (GND));
      wire XNOR_1_1_NAND5_NUM740_OUT, XNOR_1_2_NAND5_NUM740_OUT, XNOR_1_3_NAND5_NUM740_OUT;
      NOR2_X1 XNOR_1_1_NAND5_NUM740 (.ZN (XNOR_1_1_NAND5_NUM740_OUT), .A1 (N2385), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND5_NUM740 (.ZN (XNOR_1_2_NAND5_NUM740_OUT), .A1 (GND), .A2 (N2427));
      NOR2_X1 XNOR_1_3_NAND5_NUM740 (.ZN (XNOR_1_3_NAND5_NUM740_OUT), .A1 (XNOR_1_1_NAND5_NUM740_OUT), .A2 (XNOR_1_2_NAND5_NUM740_OUT));

      wire XNOR_2_1_NAND5_NUM740_OUT, XNOR_2_2_NAND5_NUM740_OUT, XNOR_2_3_NAND5_NUM740_OUT;
      NOR2_X1 XNOR_2_1_NAND5_NUM740 (.ZN (XNOR_2_1_NAND5_NUM740_OUT), .A1 (N2340), .A2 (GND));
      NOR2_X1 XNOR_2_2_NAND5_NUM740 (.ZN (XNOR_2_2_NAND5_NUM740_OUT), .A1 (GND), .A2 (N2104));
      NOR2_X1 XNOR_2_3_NAND5_NUM740 (.ZN (XNOR_2_3_NAND5_NUM740_OUT), .A1 (XNOR_2_1_NAND5_NUM740_OUT), .A2 (XNOR_2_2_NAND5_NUM740_OUT));

      wire XNOR_3_1_NAND5_NUM740_OUT, XNOR_3_2_NAND5_NUM740_OUT, XNOR_3_3_NAND5_NUM740_OUT;
      NOR2_X1 XNOR_3_1_NAND5_NUM740 (.ZN (XNOR_3_1_NAND5_NUM740_OUT), .A1 (XNOR_1_3_NAND5_NUM740_OUT), .A2 (GND));
      NOR2_X1 XNOR_3_2_NAND5_NUM740 (.ZN (XNOR_3_2_NAND5_NUM740_OUT), .A1 (GND), .A2 (XNOR_2_3_NAND5_NUM740_OUT));
      NOR2_X1 XNOR_3_3_NAND5_NUM740 (.ZN (XNOR_3_3_NAND5_NUM740_OUT), .A1 (XNOR_3_1_NAND5_NUM740_OUT), .A2 (XNOR_3_2_NAND5_NUM740_OUT));

      wire XNOR_4_1_NAND5_NUM740_OUT, XNOR_4_2_NAND5_NUM740_OUT, XNOR_4_3_NAND5_NUM740_OUT;
      NOR2_X1 XNOR_4_1_NAND5_NUM740 (.ZN (XNOR_4_1_NAND5_NUM740_OUT), .A1 (N926), .A2 (GND));
      NOR2_X1 XNOR_4_2_NAND5_NUM740 (.ZN (XNOR_4_2_NAND5_NUM740_OUT), .A1 (GND), .A2 (XNOR_3_3_NAND5_NUM740_OUT));
      NOR2_X1 XNOR_4_3_NAND5_NUM740 (.ZN (XNOR_4_3_NAND5_NUM740_OUT), .A1 (XNOR_4_1_NAND5_NUM740_OUT), .A2 (XNOR_4_2_NAND5_NUM740_OUT));

      NOR2_X1 XNOR_5_1_NAND5_NUM740 (.ZN (N2634), .A1 (XNOR_4_3_NAND5_NUM740_OUT), .A2 (GND));
      wire XNOR_1_1_AND5_NUM741_OUT, XNOR_1_2_AND5_NUM741_OUT, XNOR_1_3_AND5_NUM741_OUT;
      NOR2_X1 XNOR_1_1_AND5_NUM741 (.ZN (XNOR_1_1_AND5_NUM741_OUT), .A1 (N2286), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND5_NUM741 (.ZN (XNOR_1_2_AND5_NUM741_OUT), .A1 (GND), .A2 (N2427));
      NOR2_X1 XNOR_1_3_AND5_NUM741 (.ZN (XNOR_1_3_AND5_NUM741_OUT), .A1 (XNOR_1_1_AND5_NUM741_OUT), .A2 (XNOR_1_2_AND5_NUM741_OUT));

      wire XNOR_2_1_AND5_NUM741_OUT, XNOR_2_2_AND5_NUM741_OUT, XNOR_2_3_AND5_NUM741_OUT;
      NOR2_X1 XNOR_2_1_AND5_NUM741 (.ZN (XNOR_2_1_AND5_NUM741_OUT), .A1 (N2361), .A2 (GND));
      NOR2_X1 XNOR_2_2_AND5_NUM741 (.ZN (XNOR_2_2_AND5_NUM741_OUT), .A1 (GND), .A2 (N2129));
      NOR2_X1 XNOR_2_3_AND5_NUM741 (.ZN (XNOR_2_3_AND5_NUM741_OUT), .A1 (XNOR_2_1_AND5_NUM741_OUT), .A2 (XNOR_2_2_AND5_NUM741_OUT));

      wire XNOR_3_1_AND5_NUM741_OUT, XNOR_3_2_AND5_NUM741_OUT, XNOR_3_3_AND5_NUM741_OUT;
      NOR2_X1 XNOR_3_1_AND5_NUM741 (.ZN (XNOR_3_1_AND5_NUM741_OUT), .A1 (XNOR_1_3_AND5_NUM741_OUT), .A2 (GND));
      NOR2_X1 XNOR_3_2_AND5_NUM741 (.ZN (XNOR_3_2_AND5_NUM741_OUT), .A1 (GND), .A2 (XNOR_2_3_AND5_NUM741_OUT));
      NOR2_X1 XNOR_3_3_AND5_NUM741 (.ZN (XNOR_3_3_AND5_NUM741_OUT), .A1 (XNOR_3_1_AND5_NUM741_OUT), .A2 (XNOR_3_2_AND5_NUM741_OUT));

      wire XNOR_4_1_AND5_NUM741_OUT, XNOR_4_2_AND5_NUM741_OUT;
      NOR2_X1 XNOR_4_1_AND5_NUM741 (.ZN (XNOR_4_1_AND5_NUM741_OUT), .A1 (N1171), .A2 (GND));
      NOR2_X1 XNOR_4_2_AND5_NUM741 (.ZN (XNOR_4_2_AND5_NUM741_OUT), .A1 (GND), .A2 (XNOR_3_3_AND5_NUM741_OUT));
      NOR2_X1 XNOR_4_3_AND5_NUM741 (.ZN (N2639), .A1 (XNOR_4_1_AND5_NUM741_OUT), .A2 (XNOR_4_2_AND5_NUM741_OUT));
      wire XNOR_1_1_AND5_NUM742_OUT, XNOR_1_2_AND5_NUM742_OUT, XNOR_1_3_AND5_NUM742_OUT;
      NOR2_X1 XNOR_1_1_AND5_NUM742 (.ZN (XNOR_1_1_AND5_NUM742_OUT), .A1 (N2297), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND5_NUM742 (.ZN (XNOR_1_2_AND5_NUM742_OUT), .A1 (GND), .A2 (N2427));
      NOR2_X1 XNOR_1_3_AND5_NUM742 (.ZN (XNOR_1_3_AND5_NUM742_OUT), .A1 (XNOR_1_1_AND5_NUM742_OUT), .A2 (XNOR_1_2_AND5_NUM742_OUT));

      wire XNOR_2_1_AND5_NUM742_OUT, XNOR_2_2_AND5_NUM742_OUT, XNOR_2_3_AND5_NUM742_OUT;
      NOR2_X1 XNOR_2_1_AND5_NUM742 (.ZN (XNOR_2_1_AND5_NUM742_OUT), .A1 (N2361), .A2 (GND));
      NOR2_X1 XNOR_2_2_AND5_NUM742 (.ZN (XNOR_2_2_AND5_NUM742_OUT), .A1 (GND), .A2 (N2119));
      NOR2_X1 XNOR_2_3_AND5_NUM742 (.ZN (XNOR_2_3_AND5_NUM742_OUT), .A1 (XNOR_2_1_AND5_NUM742_OUT), .A2 (XNOR_2_2_AND5_NUM742_OUT));

      wire XNOR_3_1_AND5_NUM742_OUT, XNOR_3_2_AND5_NUM742_OUT, XNOR_3_3_AND5_NUM742_OUT;
      NOR2_X1 XNOR_3_1_AND5_NUM742 (.ZN (XNOR_3_1_AND5_NUM742_OUT), .A1 (XNOR_1_3_AND5_NUM742_OUT), .A2 (GND));
      NOR2_X1 XNOR_3_2_AND5_NUM742 (.ZN (XNOR_3_2_AND5_NUM742_OUT), .A1 (GND), .A2 (XNOR_2_3_AND5_NUM742_OUT));
      NOR2_X1 XNOR_3_3_AND5_NUM742 (.ZN (XNOR_3_3_AND5_NUM742_OUT), .A1 (XNOR_3_1_AND5_NUM742_OUT), .A2 (XNOR_3_2_AND5_NUM742_OUT));

      wire XNOR_4_1_AND5_NUM742_OUT, XNOR_4_2_AND5_NUM742_OUT;
      NOR2_X1 XNOR_4_1_AND5_NUM742 (.ZN (XNOR_4_1_AND5_NUM742_OUT), .A1 (N1171), .A2 (GND));
      NOR2_X1 XNOR_4_2_AND5_NUM742 (.ZN (XNOR_4_2_AND5_NUM742_OUT), .A1 (GND), .A2 (XNOR_3_3_AND5_NUM742_OUT));
      NOR2_X1 XNOR_4_3_AND5_NUM742 (.ZN (N2642), .A1 (XNOR_4_1_AND5_NUM742_OUT), .A2 (XNOR_4_2_AND5_NUM742_OUT));
      wire XNOR_1_1_AND5_NUM743_OUT, XNOR_1_2_AND5_NUM743_OUT, XNOR_1_3_AND5_NUM743_OUT;
      NOR2_X1 XNOR_1_1_AND5_NUM743 (.ZN (XNOR_1_1_AND5_NUM743_OUT), .A1 (N2297), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND5_NUM743 (.ZN (XNOR_1_2_AND5_NUM743_OUT), .A1 (GND), .A2 (N2427));
      NOR2_X1 XNOR_1_3_AND5_NUM743 (.ZN (XNOR_1_3_AND5_NUM743_OUT), .A1 (XNOR_1_1_AND5_NUM743_OUT), .A2 (XNOR_1_2_AND5_NUM743_OUT));

      wire XNOR_2_1_AND5_NUM743_OUT, XNOR_2_2_AND5_NUM743_OUT, XNOR_2_3_AND5_NUM743_OUT;
      NOR2_X1 XNOR_2_1_AND5_NUM743 (.ZN (XNOR_2_1_AND5_NUM743_OUT), .A1 (N2375), .A2 (GND));
      NOR2_X1 XNOR_2_2_AND5_NUM743 (.ZN (XNOR_2_2_AND5_NUM743_OUT), .A1 (GND), .A2 (N2104));
      NOR2_X1 XNOR_2_3_AND5_NUM743 (.ZN (XNOR_2_3_AND5_NUM743_OUT), .A1 (XNOR_2_1_AND5_NUM743_OUT), .A2 (XNOR_2_2_AND5_NUM743_OUT));

      wire XNOR_3_1_AND5_NUM743_OUT, XNOR_3_2_AND5_NUM743_OUT, XNOR_3_3_AND5_NUM743_OUT;
      NOR2_X1 XNOR_3_1_AND5_NUM743 (.ZN (XNOR_3_1_AND5_NUM743_OUT), .A1 (XNOR_1_3_AND5_NUM743_OUT), .A2 (GND));
      NOR2_X1 XNOR_3_2_AND5_NUM743 (.ZN (XNOR_3_2_AND5_NUM743_OUT), .A1 (GND), .A2 (XNOR_2_3_AND5_NUM743_OUT));
      NOR2_X1 XNOR_3_3_AND5_NUM743 (.ZN (XNOR_3_3_AND5_NUM743_OUT), .A1 (XNOR_3_1_AND5_NUM743_OUT), .A2 (XNOR_3_2_AND5_NUM743_OUT));

      wire XNOR_4_1_AND5_NUM743_OUT, XNOR_4_2_AND5_NUM743_OUT;
      NOR2_X1 XNOR_4_1_AND5_NUM743 (.ZN (XNOR_4_1_AND5_NUM743_OUT), .A1 (N1171), .A2 (GND));
      NOR2_X1 XNOR_4_2_AND5_NUM743 (.ZN (XNOR_4_2_AND5_NUM743_OUT), .A1 (GND), .A2 (XNOR_3_3_AND5_NUM743_OUT));
      NOR2_X1 XNOR_4_3_AND5_NUM743 (.ZN (N2645), .A1 (XNOR_4_1_AND5_NUM743_OUT), .A2 (XNOR_4_2_AND5_NUM743_OUT));
      wire XNOR_1_1_AND5_NUM744_OUT, XNOR_1_2_AND5_NUM744_OUT, XNOR_1_3_AND5_NUM744_OUT;
      NOR2_X1 XNOR_1_1_AND5_NUM744 (.ZN (XNOR_1_1_AND5_NUM744_OUT), .A1 (N2297), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND5_NUM744 (.ZN (XNOR_1_2_AND5_NUM744_OUT), .A1 (GND), .A2 (N2427));
      NOR2_X1 XNOR_1_3_AND5_NUM744 (.ZN (XNOR_1_3_AND5_NUM744_OUT), .A1 (XNOR_1_1_AND5_NUM744_OUT), .A2 (XNOR_1_2_AND5_NUM744_OUT));

      wire XNOR_2_1_AND5_NUM744_OUT, XNOR_2_2_AND5_NUM744_OUT, XNOR_2_3_AND5_NUM744_OUT;
      NOR2_X1 XNOR_2_1_AND5_NUM744 (.ZN (XNOR_2_1_AND5_NUM744_OUT), .A1 (N2340), .A2 (GND));
      NOR2_X1 XNOR_2_2_AND5_NUM744 (.ZN (XNOR_2_2_AND5_NUM744_OUT), .A1 (GND), .A2 (N2143));
      NOR2_X1 XNOR_2_3_AND5_NUM744 (.ZN (XNOR_2_3_AND5_NUM744_OUT), .A1 (XNOR_2_1_AND5_NUM744_OUT), .A2 (XNOR_2_2_AND5_NUM744_OUT));

      wire XNOR_3_1_AND5_NUM744_OUT, XNOR_3_2_AND5_NUM744_OUT, XNOR_3_3_AND5_NUM744_OUT;
      NOR2_X1 XNOR_3_1_AND5_NUM744 (.ZN (XNOR_3_1_AND5_NUM744_OUT), .A1 (XNOR_1_3_AND5_NUM744_OUT), .A2 (GND));
      NOR2_X1 XNOR_3_2_AND5_NUM744 (.ZN (XNOR_3_2_AND5_NUM744_OUT), .A1 (GND), .A2 (XNOR_2_3_AND5_NUM744_OUT));
      NOR2_X1 XNOR_3_3_AND5_NUM744 (.ZN (XNOR_3_3_AND5_NUM744_OUT), .A1 (XNOR_3_1_AND5_NUM744_OUT), .A2 (XNOR_3_2_AND5_NUM744_OUT));

      wire XNOR_4_1_AND5_NUM744_OUT, XNOR_4_2_AND5_NUM744_OUT;
      NOR2_X1 XNOR_4_1_AND5_NUM744 (.ZN (XNOR_4_1_AND5_NUM744_OUT), .A1 (N1171), .A2 (GND));
      NOR2_X1 XNOR_4_2_AND5_NUM744 (.ZN (XNOR_4_2_AND5_NUM744_OUT), .A1 (GND), .A2 (XNOR_3_3_AND5_NUM744_OUT));
      NOR2_X1 XNOR_4_3_AND5_NUM744 (.ZN (N2648), .A1 (XNOR_4_1_AND5_NUM744_OUT), .A2 (XNOR_4_2_AND5_NUM744_OUT));
      wire XNOR_1_1_AND5_NUM745_OUT, XNOR_1_2_AND5_NUM745_OUT, XNOR_1_3_AND5_NUM745_OUT;
      NOR2_X1 XNOR_1_1_AND5_NUM745 (.ZN (XNOR_1_1_AND5_NUM745_OUT), .A1 (N2297), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND5_NUM745 (.ZN (XNOR_1_2_AND5_NUM745_OUT), .A1 (GND), .A2 (N2427));
      NOR2_X1 XNOR_1_3_AND5_NUM745 (.ZN (XNOR_1_3_AND5_NUM745_OUT), .A1 (XNOR_1_1_AND5_NUM745_OUT), .A2 (XNOR_1_2_AND5_NUM745_OUT));

      wire XNOR_2_1_AND5_NUM745_OUT, XNOR_2_2_AND5_NUM745_OUT, XNOR_2_3_AND5_NUM745_OUT;
      NOR2_X1 XNOR_2_1_AND5_NUM745 (.ZN (XNOR_2_1_AND5_NUM745_OUT), .A1 (N2353), .A2 (GND));
      NOR2_X1 XNOR_2_2_AND5_NUM745 (.ZN (XNOR_2_2_AND5_NUM745_OUT), .A1 (GND), .A2 (N2129));
      NOR2_X1 XNOR_2_3_AND5_NUM745 (.ZN (XNOR_2_3_AND5_NUM745_OUT), .A1 (XNOR_2_1_AND5_NUM745_OUT), .A2 (XNOR_2_2_AND5_NUM745_OUT));

      wire XNOR_3_1_AND5_NUM745_OUT, XNOR_3_2_AND5_NUM745_OUT, XNOR_3_3_AND5_NUM745_OUT;
      NOR2_X1 XNOR_3_1_AND5_NUM745 (.ZN (XNOR_3_1_AND5_NUM745_OUT), .A1 (XNOR_1_3_AND5_NUM745_OUT), .A2 (GND));
      NOR2_X1 XNOR_3_2_AND5_NUM745 (.ZN (XNOR_3_2_AND5_NUM745_OUT), .A1 (GND), .A2 (XNOR_2_3_AND5_NUM745_OUT));
      NOR2_X1 XNOR_3_3_AND5_NUM745 (.ZN (XNOR_3_3_AND5_NUM745_OUT), .A1 (XNOR_3_1_AND5_NUM745_OUT), .A2 (XNOR_3_2_AND5_NUM745_OUT));

      wire XNOR_4_1_AND5_NUM745_OUT, XNOR_4_2_AND5_NUM745_OUT;
      NOR2_X1 XNOR_4_1_AND5_NUM745 (.ZN (XNOR_4_1_AND5_NUM745_OUT), .A1 (N1188), .A2 (GND));
      NOR2_X1 XNOR_4_2_AND5_NUM745 (.ZN (XNOR_4_2_AND5_NUM745_OUT), .A1 (GND), .A2 (XNOR_3_3_AND5_NUM745_OUT));
      NOR2_X1 XNOR_4_3_AND5_NUM745 (.ZN (N2651), .A1 (XNOR_4_1_AND5_NUM745_OUT), .A2 (XNOR_4_2_AND5_NUM745_OUT));
      wire XNOR_1_1_AND5_NUM746_OUT, XNOR_1_2_AND5_NUM746_OUT, XNOR_1_3_AND5_NUM746_OUT;
      NOR2_X1 XNOR_1_1_AND5_NUM746 (.ZN (XNOR_1_1_AND5_NUM746_OUT), .A1 (N2386), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND5_NUM746 (.ZN (XNOR_1_2_AND5_NUM746_OUT), .A1 (GND), .A2 (N2326));
      NOR2_X1 XNOR_1_3_AND5_NUM746 (.ZN (XNOR_1_3_AND5_NUM746_OUT), .A1 (XNOR_1_1_AND5_NUM746_OUT), .A2 (XNOR_1_2_AND5_NUM746_OUT));

      wire XNOR_2_1_AND5_NUM746_OUT, XNOR_2_2_AND5_NUM746_OUT, XNOR_2_3_AND5_NUM746_OUT;
      NOR2_X1 XNOR_2_1_AND5_NUM746 (.ZN (XNOR_2_1_AND5_NUM746_OUT), .A1 (N2361), .A2 (GND));
      NOR2_X1 XNOR_2_2_AND5_NUM746 (.ZN (XNOR_2_2_AND5_NUM746_OUT), .A1 (GND), .A2 (N2129));
      NOR2_X1 XNOR_2_3_AND5_NUM746 (.ZN (XNOR_2_3_AND5_NUM746_OUT), .A1 (XNOR_2_1_AND5_NUM746_OUT), .A2 (XNOR_2_2_AND5_NUM746_OUT));

      wire XNOR_3_1_AND5_NUM746_OUT, XNOR_3_2_AND5_NUM746_OUT, XNOR_3_3_AND5_NUM746_OUT;
      NOR2_X1 XNOR_3_1_AND5_NUM746 (.ZN (XNOR_3_1_AND5_NUM746_OUT), .A1 (XNOR_1_3_AND5_NUM746_OUT), .A2 (GND));
      NOR2_X1 XNOR_3_2_AND5_NUM746 (.ZN (XNOR_3_2_AND5_NUM746_OUT), .A1 (GND), .A2 (XNOR_2_3_AND5_NUM746_OUT));
      NOR2_X1 XNOR_3_3_AND5_NUM746 (.ZN (XNOR_3_3_AND5_NUM746_OUT), .A1 (XNOR_3_1_AND5_NUM746_OUT), .A2 (XNOR_3_2_AND5_NUM746_OUT));

      wire XNOR_4_1_AND5_NUM746_OUT, XNOR_4_2_AND5_NUM746_OUT;
      NOR2_X1 XNOR_4_1_AND5_NUM746 (.ZN (XNOR_4_1_AND5_NUM746_OUT), .A1 (N1188), .A2 (GND));
      NOR2_X1 XNOR_4_2_AND5_NUM746 (.ZN (XNOR_4_2_AND5_NUM746_OUT), .A1 (GND), .A2 (XNOR_3_3_AND5_NUM746_OUT));
      NOR2_X1 XNOR_4_3_AND5_NUM746 (.ZN (N2655), .A1 (XNOR_4_1_AND5_NUM746_OUT), .A2 (XNOR_4_2_AND5_NUM746_OUT));
      wire XNOR_1_1_AND5_NUM747_OUT, XNOR_1_2_AND5_NUM747_OUT, XNOR_1_3_AND5_NUM747_OUT;
      NOR2_X1 XNOR_1_1_AND5_NUM747 (.ZN (XNOR_1_1_AND5_NUM747_OUT), .A1 (N2386), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND5_NUM747 (.ZN (XNOR_1_2_AND5_NUM747_OUT), .A1 (GND), .A2 (N2326));
      NOR2_X1 XNOR_1_3_AND5_NUM747 (.ZN (XNOR_1_3_AND5_NUM747_OUT), .A1 (XNOR_1_1_AND5_NUM747_OUT), .A2 (XNOR_1_2_AND5_NUM747_OUT));

      wire XNOR_2_1_AND5_NUM747_OUT, XNOR_2_2_AND5_NUM747_OUT, XNOR_2_3_AND5_NUM747_OUT;
      NOR2_X1 XNOR_2_1_AND5_NUM747 (.ZN (XNOR_2_1_AND5_NUM747_OUT), .A1 (N2361), .A2 (GND));
      NOR2_X1 XNOR_2_2_AND5_NUM747 (.ZN (XNOR_2_2_AND5_NUM747_OUT), .A1 (GND), .A2 (N2119));
      NOR2_X1 XNOR_2_3_AND5_NUM747 (.ZN (XNOR_2_3_AND5_NUM747_OUT), .A1 (XNOR_2_1_AND5_NUM747_OUT), .A2 (XNOR_2_2_AND5_NUM747_OUT));

      wire XNOR_3_1_AND5_NUM747_OUT, XNOR_3_2_AND5_NUM747_OUT, XNOR_3_3_AND5_NUM747_OUT;
      NOR2_X1 XNOR_3_1_AND5_NUM747 (.ZN (XNOR_3_1_AND5_NUM747_OUT), .A1 (XNOR_1_3_AND5_NUM747_OUT), .A2 (GND));
      NOR2_X1 XNOR_3_2_AND5_NUM747 (.ZN (XNOR_3_2_AND5_NUM747_OUT), .A1 (GND), .A2 (XNOR_2_3_AND5_NUM747_OUT));
      NOR2_X1 XNOR_3_3_AND5_NUM747 (.ZN (XNOR_3_3_AND5_NUM747_OUT), .A1 (XNOR_3_1_AND5_NUM747_OUT), .A2 (XNOR_3_2_AND5_NUM747_OUT));

      wire XNOR_4_1_AND5_NUM747_OUT, XNOR_4_2_AND5_NUM747_OUT;
      NOR2_X1 XNOR_4_1_AND5_NUM747 (.ZN (XNOR_4_1_AND5_NUM747_OUT), .A1 (N1188), .A2 (GND));
      NOR2_X1 XNOR_4_2_AND5_NUM747 (.ZN (XNOR_4_2_AND5_NUM747_OUT), .A1 (GND), .A2 (XNOR_3_3_AND5_NUM747_OUT));
      NOR2_X1 XNOR_4_3_AND5_NUM747 (.ZN (N2658), .A1 (XNOR_4_1_AND5_NUM747_OUT), .A2 (XNOR_4_2_AND5_NUM747_OUT));
      wire XNOR_1_1_AND5_NUM748_OUT, XNOR_1_2_AND5_NUM748_OUT, XNOR_1_3_AND5_NUM748_OUT;
      NOR2_X1 XNOR_1_1_AND5_NUM748 (.ZN (XNOR_1_1_AND5_NUM748_OUT), .A1 (N2386), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND5_NUM748 (.ZN (XNOR_1_2_AND5_NUM748_OUT), .A1 (GND), .A2 (N2326));
      NOR2_X1 XNOR_1_3_AND5_NUM748 (.ZN (XNOR_1_3_AND5_NUM748_OUT), .A1 (XNOR_1_1_AND5_NUM748_OUT), .A2 (XNOR_1_2_AND5_NUM748_OUT));

      wire XNOR_2_1_AND5_NUM748_OUT, XNOR_2_2_AND5_NUM748_OUT, XNOR_2_3_AND5_NUM748_OUT;
      NOR2_X1 XNOR_2_1_AND5_NUM748 (.ZN (XNOR_2_1_AND5_NUM748_OUT), .A1 (N2375), .A2 (GND));
      NOR2_X1 XNOR_2_2_AND5_NUM748 (.ZN (XNOR_2_2_AND5_NUM748_OUT), .A1 (GND), .A2 (N2104));
      NOR2_X1 XNOR_2_3_AND5_NUM748 (.ZN (XNOR_2_3_AND5_NUM748_OUT), .A1 (XNOR_2_1_AND5_NUM748_OUT), .A2 (XNOR_2_2_AND5_NUM748_OUT));

      wire XNOR_3_1_AND5_NUM748_OUT, XNOR_3_2_AND5_NUM748_OUT, XNOR_3_3_AND5_NUM748_OUT;
      NOR2_X1 XNOR_3_1_AND5_NUM748 (.ZN (XNOR_3_1_AND5_NUM748_OUT), .A1 (XNOR_1_3_AND5_NUM748_OUT), .A2 (GND));
      NOR2_X1 XNOR_3_2_AND5_NUM748 (.ZN (XNOR_3_2_AND5_NUM748_OUT), .A1 (GND), .A2 (XNOR_2_3_AND5_NUM748_OUT));
      NOR2_X1 XNOR_3_3_AND5_NUM748 (.ZN (XNOR_3_3_AND5_NUM748_OUT), .A1 (XNOR_3_1_AND5_NUM748_OUT), .A2 (XNOR_3_2_AND5_NUM748_OUT));

      wire XNOR_4_1_AND5_NUM748_OUT, XNOR_4_2_AND5_NUM748_OUT;
      NOR2_X1 XNOR_4_1_AND5_NUM748 (.ZN (XNOR_4_1_AND5_NUM748_OUT), .A1 (N1188), .A2 (GND));
      NOR2_X1 XNOR_4_2_AND5_NUM748 (.ZN (XNOR_4_2_AND5_NUM748_OUT), .A1 (GND), .A2 (XNOR_3_3_AND5_NUM748_OUT));
      NOR2_X1 XNOR_4_3_AND5_NUM748 (.ZN (N2661), .A1 (XNOR_4_1_AND5_NUM748_OUT), .A2 (XNOR_4_2_AND5_NUM748_OUT));
      wire XNOR_1_1_AND5_NUM749_OUT, XNOR_1_2_AND5_NUM749_OUT, XNOR_1_3_AND5_NUM749_OUT;
      NOR2_X1 XNOR_1_1_AND5_NUM749 (.ZN (XNOR_1_1_AND5_NUM749_OUT), .A1 (N2386), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND5_NUM749 (.ZN (XNOR_1_2_AND5_NUM749_OUT), .A1 (GND), .A2 (N2326));
      NOR2_X1 XNOR_1_3_AND5_NUM749 (.ZN (XNOR_1_3_AND5_NUM749_OUT), .A1 (XNOR_1_1_AND5_NUM749_OUT), .A2 (XNOR_1_2_AND5_NUM749_OUT));

      wire XNOR_2_1_AND5_NUM749_OUT, XNOR_2_2_AND5_NUM749_OUT, XNOR_2_3_AND5_NUM749_OUT;
      NOR2_X1 XNOR_2_1_AND5_NUM749 (.ZN (XNOR_2_1_AND5_NUM749_OUT), .A1 (N2353), .A2 (GND));
      NOR2_X1 XNOR_2_2_AND5_NUM749 (.ZN (XNOR_2_2_AND5_NUM749_OUT), .A1 (GND), .A2 (N2129));
      NOR2_X1 XNOR_2_3_AND5_NUM749 (.ZN (XNOR_2_3_AND5_NUM749_OUT), .A1 (XNOR_2_1_AND5_NUM749_OUT), .A2 (XNOR_2_2_AND5_NUM749_OUT));

      wire XNOR_3_1_AND5_NUM749_OUT, XNOR_3_2_AND5_NUM749_OUT, XNOR_3_3_AND5_NUM749_OUT;
      NOR2_X1 XNOR_3_1_AND5_NUM749 (.ZN (XNOR_3_1_AND5_NUM749_OUT), .A1 (XNOR_1_3_AND5_NUM749_OUT), .A2 (GND));
      NOR2_X1 XNOR_3_2_AND5_NUM749 (.ZN (XNOR_3_2_AND5_NUM749_OUT), .A1 (GND), .A2 (XNOR_2_3_AND5_NUM749_OUT));
      NOR2_X1 XNOR_3_3_AND5_NUM749 (.ZN (XNOR_3_3_AND5_NUM749_OUT), .A1 (XNOR_3_1_AND5_NUM749_OUT), .A2 (XNOR_3_2_AND5_NUM749_OUT));

      wire XNOR_4_1_AND5_NUM749_OUT, XNOR_4_2_AND5_NUM749_OUT;
      NOR2_X1 XNOR_4_1_AND5_NUM749 (.ZN (XNOR_4_1_AND5_NUM749_OUT), .A1 (N1188), .A2 (GND));
      NOR2_X1 XNOR_4_2_AND5_NUM749 (.ZN (XNOR_4_2_AND5_NUM749_OUT), .A1 (GND), .A2 (XNOR_3_3_AND5_NUM749_OUT));
      NOR2_X1 XNOR_4_3_AND5_NUM749 (.ZN (N2664), .A1 (XNOR_4_1_AND5_NUM749_OUT), .A2 (XNOR_4_2_AND5_NUM749_OUT));
      wire XNOR_1_1_NAND2_NUM750_OUT, XNOR_1_2_NAND2_NUM750_OUT, XNOR_1_3_NAND2_NUM750_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM750 (.ZN (XNOR_1_1_NAND2_NUM750_OUT), .A1 (N2558), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM750 (.ZN (XNOR_1_2_NAND2_NUM750_OUT), .A1 (GND), .A2 (N534));
      NOR2_X1 XNOR_1_3_NAND2_NUM750 (.ZN (XNOR_1_3_NAND2_NUM750_OUT), .A1 (XNOR_1_1_NAND2_NUM750_OUT), .A2 (XNOR_1_2_NAND2_NUM750_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM750 (.ZN (N2669), .A1 (XNOR_1_3_NAND2_NUM750_OUT), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM751 (.ZN (N2670), .A1 (N2558), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM752_OUT, XNOR_1_2_NAND2_NUM752_OUT, XNOR_1_3_NAND2_NUM752_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM752 (.ZN (XNOR_1_1_NAND2_NUM752_OUT), .A1 (N2561), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM752 (.ZN (XNOR_1_2_NAND2_NUM752_OUT), .A1 (GND), .A2 (N535));
      NOR2_X1 XNOR_1_3_NAND2_NUM752 (.ZN (XNOR_1_3_NAND2_NUM752_OUT), .A1 (XNOR_1_1_NAND2_NUM752_OUT), .A2 (XNOR_1_2_NAND2_NUM752_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM752 (.ZN (N2671), .A1 (XNOR_1_3_NAND2_NUM752_OUT), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM753 (.ZN (N2672), .A1 (N2561), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM754_OUT, XNOR_1_2_NAND2_NUM754_OUT, XNOR_1_3_NAND2_NUM754_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM754 (.ZN (XNOR_1_1_NAND2_NUM754_OUT), .A1 (N2564), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM754 (.ZN (XNOR_1_2_NAND2_NUM754_OUT), .A1 (GND), .A2 (N536));
      NOR2_X1 XNOR_1_3_NAND2_NUM754 (.ZN (XNOR_1_3_NAND2_NUM754_OUT), .A1 (XNOR_1_1_NAND2_NUM754_OUT), .A2 (XNOR_1_2_NAND2_NUM754_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM754 (.ZN (N2673), .A1 (XNOR_1_3_NAND2_NUM754_OUT), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM755 (.ZN (N2674), .A1 (N2564), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM756_OUT, XNOR_1_2_NAND2_NUM756_OUT, XNOR_1_3_NAND2_NUM756_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM756 (.ZN (XNOR_1_1_NAND2_NUM756_OUT), .A1 (N2567), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM756 (.ZN (XNOR_1_2_NAND2_NUM756_OUT), .A1 (GND), .A2 (N537));
      NOR2_X1 XNOR_1_3_NAND2_NUM756 (.ZN (XNOR_1_3_NAND2_NUM756_OUT), .A1 (XNOR_1_1_NAND2_NUM756_OUT), .A2 (XNOR_1_2_NAND2_NUM756_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM756 (.ZN (N2675), .A1 (XNOR_1_3_NAND2_NUM756_OUT), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM757 (.ZN (N2676), .A1 (N2567), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM758_OUT, XNOR_1_2_NAND2_NUM758_OUT, XNOR_1_3_NAND2_NUM758_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM758 (.ZN (XNOR_1_1_NAND2_NUM758_OUT), .A1 (N2570), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM758 (.ZN (XNOR_1_2_NAND2_NUM758_OUT), .A1 (GND), .A2 (N543));
      NOR2_X1 XNOR_1_3_NAND2_NUM758 (.ZN (XNOR_1_3_NAND2_NUM758_OUT), .A1 (XNOR_1_1_NAND2_NUM758_OUT), .A2 (XNOR_1_2_NAND2_NUM758_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM758 (.ZN (N2682), .A1 (XNOR_1_3_NAND2_NUM758_OUT), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM759 (.ZN (N2683), .A1 (N2570), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM760_OUT, XNOR_1_2_NAND2_NUM760_OUT, XNOR_1_3_NAND2_NUM760_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM760 (.ZN (XNOR_1_1_NAND2_NUM760_OUT), .A1 (N2573), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM760 (.ZN (XNOR_1_2_NAND2_NUM760_OUT), .A1 (GND), .A2 (N548));
      NOR2_X1 XNOR_1_3_NAND2_NUM760 (.ZN (XNOR_1_3_NAND2_NUM760_OUT), .A1 (XNOR_1_1_NAND2_NUM760_OUT), .A2 (XNOR_1_2_NAND2_NUM760_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM760 (.ZN (N2688), .A1 (XNOR_1_3_NAND2_NUM760_OUT), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM761 (.ZN (N2689), .A1 (N2573), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM762_OUT, XNOR_1_2_NAND2_NUM762_OUT, XNOR_1_3_NAND2_NUM762_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM762 (.ZN (XNOR_1_1_NAND2_NUM762_OUT), .A1 (N2576), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM762 (.ZN (XNOR_1_2_NAND2_NUM762_OUT), .A1 (GND), .A2 (N549));
      NOR2_X1 XNOR_1_3_NAND2_NUM762 (.ZN (XNOR_1_3_NAND2_NUM762_OUT), .A1 (XNOR_1_1_NAND2_NUM762_OUT), .A2 (XNOR_1_2_NAND2_NUM762_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM762 (.ZN (N2690), .A1 (XNOR_1_3_NAND2_NUM762_OUT), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM763 (.ZN (N2691), .A1 (N2576), .A2 (GND));
      wire XNOR_1_1_AND8_NUM764_OUT, XNOR_1_2_AND8_NUM764_OUT, XNOR_1_3_AND8_NUM764_OUT;
      NOR2_X1 XNOR_1_1_AND8_NUM764 (.ZN (XNOR_1_1_AND8_NUM764_OUT), .A1 (N2627), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND8_NUM764 (.ZN (XNOR_1_2_AND8_NUM764_OUT), .A1 (GND), .A2 (N2628));
      NOR2_X1 XNOR_1_3_AND8_NUM764 (.ZN (XNOR_1_3_AND8_NUM764_OUT), .A1 (XNOR_1_1_AND8_NUM764_OUT), .A2 (XNOR_1_2_AND8_NUM764_OUT));

      wire XNOR_2_1_AND8_NUM764_OUT, XNOR_2_2_AND8_NUM764_OUT, XNOR_2_3_AND8_NUM764_OUT;
      NOR2_X1 XNOR_2_1_AND8_NUM764 (.ZN (XNOR_2_1_AND8_NUM764_OUT), .A1 (N2629), .A2 (GND));
      NOR2_X1 XNOR_2_2_AND8_NUM764 (.ZN (XNOR_2_2_AND8_NUM764_OUT), .A1 (GND), .A2 (N2630));
      NOR2_X1 XNOR_2_3_AND8_NUM764 (.ZN (XNOR_2_3_AND8_NUM764_OUT), .A1 (XNOR_2_1_AND8_NUM764_OUT), .A2 (XNOR_2_2_AND8_NUM764_OUT));

      wire XNOR_3_1_AND8_NUM764_OUT, XNOR_3_2_AND8_NUM764_OUT, XNOR_3_3_AND8_NUM764_OUT;
      NOR2_X1 XNOR_3_1_AND8_NUM764 (.ZN (XNOR_3_1_AND8_NUM764_OUT), .A1 (N2631), .A2 (GND));
      NOR2_X1 XNOR_3_2_AND8_NUM764 (.ZN (XNOR_3_2_AND8_NUM764_OUT), .A1 (GND), .A2 (N2632));
      NOR2_X1 XNOR_3_3_AND8_NUM764 (.ZN (XNOR_3_3_AND8_NUM764_OUT), .A1 (XNOR_3_1_AND8_NUM764_OUT), .A2 (XNOR_3_2_AND8_NUM764_OUT));

      wire XNOR_4_1_AND8_NUM764_OUT, XNOR_4_2_AND8_NUM764_OUT, XNOR_4_3_AND8_NUM764_OUT;
      NOR2_X1 XNOR_4_1_AND8_NUM764 (.ZN (XNOR_4_1_AND8_NUM764_OUT), .A1 (N2633), .A2 (GND));
      NOR2_X1 XNOR_4_2_AND8_NUM764 (.ZN (XNOR_4_2_AND8_NUM764_OUT), .A1 (GND), .A2 (N2634));
      NOR2_X1 XNOR_4_3_AND8_NUM764 (.ZN (XNOR_4_3_AND8_NUM764_OUT), .A1 (XNOR_4_1_AND8_NUM764_OUT), .A2 (XNOR_4_2_AND8_NUM764_OUT));

      wire XNOR_5_1_AND8_NUM764_OUT, XNOR_5_2_AND8_NUM764_OUT, XNOR_5_3_AND8_NUM764_OUT;
      NOR2_X1 XNOR_5_1_AND8_NUM764 (.ZN (XNOR_5_1_AND8_NUM764_OUT), .A1 (XNOR_1_3_AND8_NUM764_OUT), .A2 (GND));
      NOR2_X1 XNOR_5_2_AND8_NUM764 (.ZN (XNOR_5_2_AND8_NUM764_OUT), .A1 (GND), .A2 (XNOR_2_3_AND8_NUM764_OUT));
      NOR2_X1 XNOR_5_3_AND8_NUM764 (.ZN (XNOR_5_3_AND8_NUM764_OUT), .A1 (XNOR_5_1_AND8_NUM764_OUT), .A2 (XNOR_5_2_AND8_NUM764_OUT));

      wire XNOR_6_1_AND8_NUM764_OUT, XNOR_6_2_AND8_NUM764_OUT, XNOR_6_3_AND8_NUM764_OUT;
      NOR2_X1 XNOR_6_1_AND8_NUM764 (.ZN (XNOR_6_1_AND8_NUM764_OUT), .A1 (XNOR_3_3_AND8_NUM764_OUT), .A2 (GND));
      NOR2_X1 XNOR_6_2_AND8_NUM764 (.ZN (XNOR_6_2_AND8_NUM764_OUT), .A1 (GND), .A2 (XNOR_4_3_AND8_NUM764_OUT));
      NOR2_X1 XNOR_6_3_AND8_NUM764 (.ZN (XNOR_6_3_AND8_NUM764_OUT), .A1 (XNOR_6_1_AND8_NUM764_OUT), .A2 (XNOR_6_2_AND8_NUM764_OUT));

      wire XNOR_7_1_AND8_NUM764_OUT, XNOR_7_2_AND8_NUM764_OUT;
      NOR2_X1 XNOR_7_1_AND8_NUM764 (.ZN (XNOR_7_1_AND8_NUM764_OUT), .A1 (XNOR_5_3_AND8_NUM764_OUT), .A2 (GND));
      NOR2_X1 XNOR_7_2_AND8_NUM764 (.ZN (XNOR_7_2_AND8_NUM764_OUT), .A1 (GND), .A2 (XNOR_6_3_AND8_NUM764_OUT));
      NOR2_X1 XNOR_7_3_AND8_NUM764 (.ZN (N2710), .A1 (XNOR_7_1_AND8_NUM764_OUT), .A2 (XNOR_7_2_AND8_NUM764_OUT));
      wire XNOR_1_1_NAND2_NUM765_OUT, XNOR_1_2_NAND2_NUM765_OUT, XNOR_1_3_NAND2_NUM765_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM765 (.ZN (XNOR_1_1_NAND2_NUM765_OUT), .A1 (N343), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM765 (.ZN (XNOR_1_2_NAND2_NUM765_OUT), .A1 (GND), .A2 (N2670));
      NOR2_X1 XNOR_1_3_NAND2_NUM765 (.ZN (XNOR_1_3_NAND2_NUM765_OUT), .A1 (XNOR_1_1_NAND2_NUM765_OUT), .A2 (XNOR_1_2_NAND2_NUM765_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM765 (.ZN (N2720), .A1 (XNOR_1_3_NAND2_NUM765_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM766_OUT, XNOR_1_2_NAND2_NUM766_OUT, XNOR_1_3_NAND2_NUM766_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM766 (.ZN (XNOR_1_1_NAND2_NUM766_OUT), .A1 (N346), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM766 (.ZN (XNOR_1_2_NAND2_NUM766_OUT), .A1 (GND), .A2 (N2672));
      NOR2_X1 XNOR_1_3_NAND2_NUM766 (.ZN (XNOR_1_3_NAND2_NUM766_OUT), .A1 (XNOR_1_1_NAND2_NUM766_OUT), .A2 (XNOR_1_2_NAND2_NUM766_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM766 (.ZN (N2721), .A1 (XNOR_1_3_NAND2_NUM766_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM767_OUT, XNOR_1_2_NAND2_NUM767_OUT, XNOR_1_3_NAND2_NUM767_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM767 (.ZN (XNOR_1_1_NAND2_NUM767_OUT), .A1 (N349), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM767 (.ZN (XNOR_1_2_NAND2_NUM767_OUT), .A1 (GND), .A2 (N2674));
      NOR2_X1 XNOR_1_3_NAND2_NUM767 (.ZN (XNOR_1_3_NAND2_NUM767_OUT), .A1 (XNOR_1_1_NAND2_NUM767_OUT), .A2 (XNOR_1_2_NAND2_NUM767_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM767 (.ZN (N2722), .A1 (XNOR_1_3_NAND2_NUM767_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM768_OUT, XNOR_1_2_NAND2_NUM768_OUT, XNOR_1_3_NAND2_NUM768_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM768 (.ZN (XNOR_1_1_NAND2_NUM768_OUT), .A1 (N352), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM768 (.ZN (XNOR_1_2_NAND2_NUM768_OUT), .A1 (GND), .A2 (N2676));
      NOR2_X1 XNOR_1_3_NAND2_NUM768 (.ZN (XNOR_1_3_NAND2_NUM768_OUT), .A1 (XNOR_1_1_NAND2_NUM768_OUT), .A2 (XNOR_1_2_NAND2_NUM768_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM768 (.ZN (N2723), .A1 (XNOR_1_3_NAND2_NUM768_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM769_OUT, XNOR_1_2_NAND2_NUM769_OUT, XNOR_1_3_NAND2_NUM769_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM769 (.ZN (XNOR_1_1_NAND2_NUM769_OUT), .A1 (N2639), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM769 (.ZN (XNOR_1_2_NAND2_NUM769_OUT), .A1 (GND), .A2 (N538));
      NOR2_X1 XNOR_1_3_NAND2_NUM769 (.ZN (XNOR_1_3_NAND2_NUM769_OUT), .A1 (XNOR_1_1_NAND2_NUM769_OUT), .A2 (XNOR_1_2_NAND2_NUM769_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM769 (.ZN (N2724), .A1 (XNOR_1_3_NAND2_NUM769_OUT), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM770 (.ZN (N2725), .A1 (N2639), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM771_OUT, XNOR_1_2_NAND2_NUM771_OUT, XNOR_1_3_NAND2_NUM771_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM771 (.ZN (XNOR_1_1_NAND2_NUM771_OUT), .A1 (N2642), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM771 (.ZN (XNOR_1_2_NAND2_NUM771_OUT), .A1 (GND), .A2 (N539));
      NOR2_X1 XNOR_1_3_NAND2_NUM771 (.ZN (XNOR_1_3_NAND2_NUM771_OUT), .A1 (XNOR_1_1_NAND2_NUM771_OUT), .A2 (XNOR_1_2_NAND2_NUM771_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM771 (.ZN (N2726), .A1 (XNOR_1_3_NAND2_NUM771_OUT), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM772 (.ZN (N2727), .A1 (N2642), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM773_OUT, XNOR_1_2_NAND2_NUM773_OUT, XNOR_1_3_NAND2_NUM773_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM773 (.ZN (XNOR_1_1_NAND2_NUM773_OUT), .A1 (N2645), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM773 (.ZN (XNOR_1_2_NAND2_NUM773_OUT), .A1 (GND), .A2 (N540));
      NOR2_X1 XNOR_1_3_NAND2_NUM773 (.ZN (XNOR_1_3_NAND2_NUM773_OUT), .A1 (XNOR_1_1_NAND2_NUM773_OUT), .A2 (XNOR_1_2_NAND2_NUM773_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM773 (.ZN (N2728), .A1 (XNOR_1_3_NAND2_NUM773_OUT), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM774 (.ZN (N2729), .A1 (N2645), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM775_OUT, XNOR_1_2_NAND2_NUM775_OUT, XNOR_1_3_NAND2_NUM775_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM775 (.ZN (XNOR_1_1_NAND2_NUM775_OUT), .A1 (N2648), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM775 (.ZN (XNOR_1_2_NAND2_NUM775_OUT), .A1 (GND), .A2 (N541));
      NOR2_X1 XNOR_1_3_NAND2_NUM775 (.ZN (XNOR_1_3_NAND2_NUM775_OUT), .A1 (XNOR_1_1_NAND2_NUM775_OUT), .A2 (XNOR_1_2_NAND2_NUM775_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM775 (.ZN (N2730), .A1 (XNOR_1_3_NAND2_NUM775_OUT), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM776 (.ZN (N2731), .A1 (N2648), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM777_OUT, XNOR_1_2_NAND2_NUM777_OUT, XNOR_1_3_NAND2_NUM777_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM777 (.ZN (XNOR_1_1_NAND2_NUM777_OUT), .A1 (N2651), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM777 (.ZN (XNOR_1_2_NAND2_NUM777_OUT), .A1 (GND), .A2 (N542));
      NOR2_X1 XNOR_1_3_NAND2_NUM777 (.ZN (XNOR_1_3_NAND2_NUM777_OUT), .A1 (XNOR_1_1_NAND2_NUM777_OUT), .A2 (XNOR_1_2_NAND2_NUM777_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM777 (.ZN (N2732), .A1 (XNOR_1_3_NAND2_NUM777_OUT), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM778 (.ZN (N2733), .A1 (N2651), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM779_OUT, XNOR_1_2_NAND2_NUM779_OUT, XNOR_1_3_NAND2_NUM779_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM779 (.ZN (XNOR_1_1_NAND2_NUM779_OUT), .A1 (N370), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM779 (.ZN (XNOR_1_2_NAND2_NUM779_OUT), .A1 (GND), .A2 (N2683));
      NOR2_X1 XNOR_1_3_NAND2_NUM779 (.ZN (XNOR_1_3_NAND2_NUM779_OUT), .A1 (XNOR_1_1_NAND2_NUM779_OUT), .A2 (XNOR_1_2_NAND2_NUM779_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM779 (.ZN (N2734), .A1 (XNOR_1_3_NAND2_NUM779_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM780_OUT, XNOR_1_2_NAND2_NUM780_OUT, XNOR_1_3_NAND2_NUM780_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM780 (.ZN (XNOR_1_1_NAND2_NUM780_OUT), .A1 (N2655), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM780 (.ZN (XNOR_1_2_NAND2_NUM780_OUT), .A1 (GND), .A2 (N544));
      NOR2_X1 XNOR_1_3_NAND2_NUM780 (.ZN (XNOR_1_3_NAND2_NUM780_OUT), .A1 (XNOR_1_1_NAND2_NUM780_OUT), .A2 (XNOR_1_2_NAND2_NUM780_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM780 (.ZN (N2735), .A1 (XNOR_1_3_NAND2_NUM780_OUT), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM781 (.ZN (N2736), .A1 (N2655), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM782_OUT, XNOR_1_2_NAND2_NUM782_OUT, XNOR_1_3_NAND2_NUM782_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM782 (.ZN (XNOR_1_1_NAND2_NUM782_OUT), .A1 (N2658), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM782 (.ZN (XNOR_1_2_NAND2_NUM782_OUT), .A1 (GND), .A2 (N545));
      NOR2_X1 XNOR_1_3_NAND2_NUM782 (.ZN (XNOR_1_3_NAND2_NUM782_OUT), .A1 (XNOR_1_1_NAND2_NUM782_OUT), .A2 (XNOR_1_2_NAND2_NUM782_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM782 (.ZN (N2737), .A1 (XNOR_1_3_NAND2_NUM782_OUT), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM783 (.ZN (N2738), .A1 (N2658), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM784_OUT, XNOR_1_2_NAND2_NUM784_OUT, XNOR_1_3_NAND2_NUM784_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM784 (.ZN (XNOR_1_1_NAND2_NUM784_OUT), .A1 (N2661), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM784 (.ZN (XNOR_1_2_NAND2_NUM784_OUT), .A1 (GND), .A2 (N546));
      NOR2_X1 XNOR_1_3_NAND2_NUM784 (.ZN (XNOR_1_3_NAND2_NUM784_OUT), .A1 (XNOR_1_1_NAND2_NUM784_OUT), .A2 (XNOR_1_2_NAND2_NUM784_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM784 (.ZN (N2739), .A1 (XNOR_1_3_NAND2_NUM784_OUT), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM785 (.ZN (N2740), .A1 (N2661), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM786_OUT, XNOR_1_2_NAND2_NUM786_OUT, XNOR_1_3_NAND2_NUM786_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM786 (.ZN (XNOR_1_1_NAND2_NUM786_OUT), .A1 (N2664), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM786 (.ZN (XNOR_1_2_NAND2_NUM786_OUT), .A1 (GND), .A2 (N547));
      NOR2_X1 XNOR_1_3_NAND2_NUM786 (.ZN (XNOR_1_3_NAND2_NUM786_OUT), .A1 (XNOR_1_1_NAND2_NUM786_OUT), .A2 (XNOR_1_2_NAND2_NUM786_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM786 (.ZN (N2741), .A1 (XNOR_1_3_NAND2_NUM786_OUT), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM787 (.ZN (N2742), .A1 (N2664), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM788_OUT, XNOR_1_2_NAND2_NUM788_OUT, XNOR_1_3_NAND2_NUM788_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM788 (.ZN (XNOR_1_1_NAND2_NUM788_OUT), .A1 (N385), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM788 (.ZN (XNOR_1_2_NAND2_NUM788_OUT), .A1 (GND), .A2 (N2689));
      NOR2_X1 XNOR_1_3_NAND2_NUM788 (.ZN (XNOR_1_3_NAND2_NUM788_OUT), .A1 (XNOR_1_1_NAND2_NUM788_OUT), .A2 (XNOR_1_2_NAND2_NUM788_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM788 (.ZN (N2743), .A1 (XNOR_1_3_NAND2_NUM788_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM789_OUT, XNOR_1_2_NAND2_NUM789_OUT, XNOR_1_3_NAND2_NUM789_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM789 (.ZN (XNOR_1_1_NAND2_NUM789_OUT), .A1 (N388), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM789 (.ZN (XNOR_1_2_NAND2_NUM789_OUT), .A1 (GND), .A2 (N2691));
      NOR2_X1 XNOR_1_3_NAND2_NUM789 (.ZN (XNOR_1_3_NAND2_NUM789_OUT), .A1 (XNOR_1_1_NAND2_NUM789_OUT), .A2 (XNOR_1_2_NAND2_NUM789_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM789 (.ZN (N2744), .A1 (XNOR_1_3_NAND2_NUM789_OUT), .A2 (GND));
      wire XNOR_1_1_NAND8_NUM790_OUT, XNOR_1_2_NAND8_NUM790_OUT, XNOR_1_3_NAND8_NUM790_OUT;
      NOR2_X1 XNOR_1_1_NAND8_NUM790 (.ZN (XNOR_1_1_NAND8_NUM790_OUT), .A1 (N2537), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND8_NUM790 (.ZN (XNOR_1_2_NAND8_NUM790_OUT), .A1 (GND), .A2 (N2540));
      NOR2_X1 XNOR_1_3_NAND8_NUM790 (.ZN (XNOR_1_3_NAND8_NUM790_OUT), .A1 (XNOR_1_1_NAND8_NUM790_OUT), .A2 (XNOR_1_2_NAND8_NUM790_OUT));

      wire XNOR_2_1_NAND8_NUM790_OUT, XNOR_2_2_NAND8_NUM790_OUT, XNOR_2_3_NAND8_NUM790_OUT;
      NOR2_X1 XNOR_2_1_NAND8_NUM790 (.ZN (XNOR_2_1_NAND8_NUM790_OUT), .A1 (N2543), .A2 (GND));
      NOR2_X1 XNOR_2_2_NAND8_NUM790 (.ZN (XNOR_2_2_NAND8_NUM790_OUT), .A1 (GND), .A2 (N2546));
      NOR2_X1 XNOR_2_3_NAND8_NUM790 (.ZN (XNOR_2_3_NAND8_NUM790_OUT), .A1 (XNOR_2_1_NAND8_NUM790_OUT), .A2 (XNOR_2_2_NAND8_NUM790_OUT));

      wire XNOR_3_1_NAND8_NUM790_OUT, XNOR_3_2_NAND8_NUM790_OUT, XNOR_3_3_NAND8_NUM790_OUT;
      NOR2_X1 XNOR_3_1_NAND8_NUM790 (.ZN (XNOR_3_1_NAND8_NUM790_OUT), .A1 (N2594), .A2 (GND));
      NOR2_X1 XNOR_3_2_NAND8_NUM790 (.ZN (XNOR_3_2_NAND8_NUM790_OUT), .A1 (GND), .A2 (N2597));
      NOR2_X1 XNOR_3_3_NAND8_NUM790 (.ZN (XNOR_3_3_NAND8_NUM790_OUT), .A1 (XNOR_3_1_NAND8_NUM790_OUT), .A2 (XNOR_3_2_NAND8_NUM790_OUT));

      wire XNOR_4_1_NAND8_NUM790_OUT, XNOR_4_2_NAND8_NUM790_OUT, XNOR_4_3_NAND8_NUM790_OUT;
      NOR2_X1 XNOR_4_1_NAND8_NUM790 (.ZN (XNOR_4_1_NAND8_NUM790_OUT), .A1 (N2600), .A2 (GND));
      NOR2_X1 XNOR_4_2_NAND8_NUM790 (.ZN (XNOR_4_2_NAND8_NUM790_OUT), .A1 (GND), .A2 (N2603));
      NOR2_X1 XNOR_4_3_NAND8_NUM790 (.ZN (XNOR_4_3_NAND8_NUM790_OUT), .A1 (XNOR_4_1_NAND8_NUM790_OUT), .A2 (XNOR_4_2_NAND8_NUM790_OUT));

      wire XNOR_5_1_NAND8_NUM790_OUT, XNOR_5_2_NAND8_NUM790_OUT, XNOR_5_3_NAND8_NUM790_OUT;
      NOR2_X1 XNOR_5_1_NAND8_NUM790 (.ZN (XNOR_5_1_NAND8_NUM790_OUT), .A1 (XNOR_1_3_NAND8_NUM790_OUT), .A2 (GND));
      NOR2_X1 XNOR_5_2_NAND8_NUM790 (.ZN (XNOR_5_2_NAND8_NUM790_OUT), .A1 (GND), .A2 (XNOR_2_3_NAND8_NUM790_OUT));
      NOR2_X1 XNOR_5_3_NAND8_NUM790 (.ZN (XNOR_5_3_NAND8_NUM790_OUT), .A1 (XNOR_5_1_NAND8_NUM790_OUT), .A2 (XNOR_5_2_NAND8_NUM790_OUT));

      wire XNOR_6_1_NAND8_NUM790_OUT, XNOR_6_2_NAND8_NUM790_OUT, XNOR_6_3_NAND8_NUM790_OUT;
      NOR2_X1 XNOR_6_1_NAND8_NUM790 (.ZN (XNOR_6_1_NAND8_NUM790_OUT), .A1 (XNOR_3_3_NAND8_NUM790_OUT), .A2 (GND));
      NOR2_X1 XNOR_6_2_NAND8_NUM790 (.ZN (XNOR_6_2_NAND8_NUM790_OUT), .A1 (GND), .A2 (XNOR_4_3_NAND8_NUM790_OUT));
      NOR2_X1 XNOR_6_3_NAND8_NUM790 (.ZN (XNOR_6_3_NAND8_NUM790_OUT), .A1 (XNOR_6_1_NAND8_NUM790_OUT), .A2 (XNOR_6_2_NAND8_NUM790_OUT));

      wire XNOR_7_1_NAND8_NUM790_OUT, XNOR_7_2_NAND8_NUM790_OUT, XNOR_7_3_NAND8_NUM790_OUT;
      NOR2_X1 XNOR_7_1_NAND8_NUM790 (.ZN (XNOR_7_1_NAND8_NUM790_OUT), .A1 (XNOR_5_3_NAND8_NUM790_OUT), .A2 (GND));
      NOR2_X1 XNOR_7_2_NAND8_NUM790 (.ZN (XNOR_7_2_NAND8_NUM790_OUT), .A1 (GND), .A2 (XNOR_6_3_NAND8_NUM790_OUT));
      NOR2_X1 XNOR_7_3_NAND8_NUM790 (.ZN (XNOR_7_3_NAND8_NUM790_OUT), .A1 (XNOR_7_1_NAND8_NUM790_OUT), .A2 (XNOR_7_2_NAND8_NUM790_OUT));

      NOR2_X1 XNOR_8_1_NAND8_NUM790 (.ZN (N2745), .A1 (XNOR_7_3_NAND8_NUM790_OUT), .A2 (GND));
      wire XNOR_1_1_NAND8_NUM791_OUT, XNOR_1_2_NAND8_NUM791_OUT, XNOR_1_3_NAND8_NUM791_OUT;
      NOR2_X1 XNOR_1_1_NAND8_NUM791 (.ZN (XNOR_1_1_NAND8_NUM791_OUT), .A1 (N2606), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND8_NUM791 (.ZN (XNOR_1_2_NAND8_NUM791_OUT), .A1 (GND), .A2 (N2549));
      NOR2_X1 XNOR_1_3_NAND8_NUM791 (.ZN (XNOR_1_3_NAND8_NUM791_OUT), .A1 (XNOR_1_1_NAND8_NUM791_OUT), .A2 (XNOR_1_2_NAND8_NUM791_OUT));

      wire XNOR_2_1_NAND8_NUM791_OUT, XNOR_2_2_NAND8_NUM791_OUT, XNOR_2_3_NAND8_NUM791_OUT;
      NOR2_X1 XNOR_2_1_NAND8_NUM791 (.ZN (XNOR_2_1_NAND8_NUM791_OUT), .A1 (N2611), .A2 (GND));
      NOR2_X1 XNOR_2_2_NAND8_NUM791 (.ZN (XNOR_2_2_NAND8_NUM791_OUT), .A1 (GND), .A2 (N2614));
      NOR2_X1 XNOR_2_3_NAND8_NUM791 (.ZN (XNOR_2_3_NAND8_NUM791_OUT), .A1 (XNOR_2_1_NAND8_NUM791_OUT), .A2 (XNOR_2_2_NAND8_NUM791_OUT));

      wire XNOR_3_1_NAND8_NUM791_OUT, XNOR_3_2_NAND8_NUM791_OUT, XNOR_3_3_NAND8_NUM791_OUT;
      NOR2_X1 XNOR_3_1_NAND8_NUM791 (.ZN (XNOR_3_1_NAND8_NUM791_OUT), .A1 (N2617), .A2 (GND));
      NOR2_X1 XNOR_3_2_NAND8_NUM791 (.ZN (XNOR_3_2_NAND8_NUM791_OUT), .A1 (GND), .A2 (N2620));
      NOR2_X1 XNOR_3_3_NAND8_NUM791 (.ZN (XNOR_3_3_NAND8_NUM791_OUT), .A1 (XNOR_3_1_NAND8_NUM791_OUT), .A2 (XNOR_3_2_NAND8_NUM791_OUT));

      wire XNOR_4_1_NAND8_NUM791_OUT, XNOR_4_2_NAND8_NUM791_OUT, XNOR_4_3_NAND8_NUM791_OUT;
      NOR2_X1 XNOR_4_1_NAND8_NUM791 (.ZN (XNOR_4_1_NAND8_NUM791_OUT), .A1 (N2552), .A2 (GND));
      NOR2_X1 XNOR_4_2_NAND8_NUM791 (.ZN (XNOR_4_2_NAND8_NUM791_OUT), .A1 (GND), .A2 (N2555));
      NOR2_X1 XNOR_4_3_NAND8_NUM791 (.ZN (XNOR_4_3_NAND8_NUM791_OUT), .A1 (XNOR_4_1_NAND8_NUM791_OUT), .A2 (XNOR_4_2_NAND8_NUM791_OUT));

      wire XNOR_5_1_NAND8_NUM791_OUT, XNOR_5_2_NAND8_NUM791_OUT, XNOR_5_3_NAND8_NUM791_OUT;
      NOR2_X1 XNOR_5_1_NAND8_NUM791 (.ZN (XNOR_5_1_NAND8_NUM791_OUT), .A1 (XNOR_1_3_NAND8_NUM791_OUT), .A2 (GND));
      NOR2_X1 XNOR_5_2_NAND8_NUM791 (.ZN (XNOR_5_2_NAND8_NUM791_OUT), .A1 (GND), .A2 (XNOR_2_3_NAND8_NUM791_OUT));
      NOR2_X1 XNOR_5_3_NAND8_NUM791 (.ZN (XNOR_5_3_NAND8_NUM791_OUT), .A1 (XNOR_5_1_NAND8_NUM791_OUT), .A2 (XNOR_5_2_NAND8_NUM791_OUT));

      wire XNOR_6_1_NAND8_NUM791_OUT, XNOR_6_2_NAND8_NUM791_OUT, XNOR_6_3_NAND8_NUM791_OUT;
      NOR2_X1 XNOR_6_1_NAND8_NUM791 (.ZN (XNOR_6_1_NAND8_NUM791_OUT), .A1 (XNOR_3_3_NAND8_NUM791_OUT), .A2 (GND));
      NOR2_X1 XNOR_6_2_NAND8_NUM791 (.ZN (XNOR_6_2_NAND8_NUM791_OUT), .A1 (GND), .A2 (XNOR_4_3_NAND8_NUM791_OUT));
      NOR2_X1 XNOR_6_3_NAND8_NUM791 (.ZN (XNOR_6_3_NAND8_NUM791_OUT), .A1 (XNOR_6_1_NAND8_NUM791_OUT), .A2 (XNOR_6_2_NAND8_NUM791_OUT));

      wire XNOR_7_1_NAND8_NUM791_OUT, XNOR_7_2_NAND8_NUM791_OUT, XNOR_7_3_NAND8_NUM791_OUT;
      NOR2_X1 XNOR_7_1_NAND8_NUM791 (.ZN (XNOR_7_1_NAND8_NUM791_OUT), .A1 (XNOR_5_3_NAND8_NUM791_OUT), .A2 (GND));
      NOR2_X1 XNOR_7_2_NAND8_NUM791 (.ZN (XNOR_7_2_NAND8_NUM791_OUT), .A1 (GND), .A2 (XNOR_6_3_NAND8_NUM791_OUT));
      NOR2_X1 XNOR_7_3_NAND8_NUM791 (.ZN (XNOR_7_3_NAND8_NUM791_OUT), .A1 (XNOR_7_1_NAND8_NUM791_OUT), .A2 (XNOR_7_2_NAND8_NUM791_OUT));

      NOR2_X1 XNOR_8_1_NAND8_NUM791 (.ZN (N2746), .A1 (XNOR_7_3_NAND8_NUM791_OUT), .A2 (GND));
      wire XNOR_1_1_AND8_NUM792_OUT, XNOR_1_2_AND8_NUM792_OUT, XNOR_1_3_AND8_NUM792_OUT;
      NOR2_X1 XNOR_1_1_AND8_NUM792 (.ZN (XNOR_1_1_AND8_NUM792_OUT), .A1 (N2537), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND8_NUM792 (.ZN (XNOR_1_2_AND8_NUM792_OUT), .A1 (GND), .A2 (N2540));
      NOR2_X1 XNOR_1_3_AND8_NUM792 (.ZN (XNOR_1_3_AND8_NUM792_OUT), .A1 (XNOR_1_1_AND8_NUM792_OUT), .A2 (XNOR_1_2_AND8_NUM792_OUT));

      wire XNOR_2_1_AND8_NUM792_OUT, XNOR_2_2_AND8_NUM792_OUT, XNOR_2_3_AND8_NUM792_OUT;
      NOR2_X1 XNOR_2_1_AND8_NUM792 (.ZN (XNOR_2_1_AND8_NUM792_OUT), .A1 (N2543), .A2 (GND));
      NOR2_X1 XNOR_2_2_AND8_NUM792 (.ZN (XNOR_2_2_AND8_NUM792_OUT), .A1 (GND), .A2 (N2546));
      NOR2_X1 XNOR_2_3_AND8_NUM792 (.ZN (XNOR_2_3_AND8_NUM792_OUT), .A1 (XNOR_2_1_AND8_NUM792_OUT), .A2 (XNOR_2_2_AND8_NUM792_OUT));

      wire XNOR_3_1_AND8_NUM792_OUT, XNOR_3_2_AND8_NUM792_OUT, XNOR_3_3_AND8_NUM792_OUT;
      NOR2_X1 XNOR_3_1_AND8_NUM792 (.ZN (XNOR_3_1_AND8_NUM792_OUT), .A1 (N2594), .A2 (GND));
      NOR2_X1 XNOR_3_2_AND8_NUM792 (.ZN (XNOR_3_2_AND8_NUM792_OUT), .A1 (GND), .A2 (N2597));
      NOR2_X1 XNOR_3_3_AND8_NUM792 (.ZN (XNOR_3_3_AND8_NUM792_OUT), .A1 (XNOR_3_1_AND8_NUM792_OUT), .A2 (XNOR_3_2_AND8_NUM792_OUT));

      wire XNOR_4_1_AND8_NUM792_OUT, XNOR_4_2_AND8_NUM792_OUT, XNOR_4_3_AND8_NUM792_OUT;
      NOR2_X1 XNOR_4_1_AND8_NUM792 (.ZN (XNOR_4_1_AND8_NUM792_OUT), .A1 (N2600), .A2 (GND));
      NOR2_X1 XNOR_4_2_AND8_NUM792 (.ZN (XNOR_4_2_AND8_NUM792_OUT), .A1 (GND), .A2 (N2603));
      NOR2_X1 XNOR_4_3_AND8_NUM792 (.ZN (XNOR_4_3_AND8_NUM792_OUT), .A1 (XNOR_4_1_AND8_NUM792_OUT), .A2 (XNOR_4_2_AND8_NUM792_OUT));

      wire XNOR_5_1_AND8_NUM792_OUT, XNOR_5_2_AND8_NUM792_OUT, XNOR_5_3_AND8_NUM792_OUT;
      NOR2_X1 XNOR_5_1_AND8_NUM792 (.ZN (XNOR_5_1_AND8_NUM792_OUT), .A1 (XNOR_1_3_AND8_NUM792_OUT), .A2 (GND));
      NOR2_X1 XNOR_5_2_AND8_NUM792 (.ZN (XNOR_5_2_AND8_NUM792_OUT), .A1 (GND), .A2 (XNOR_2_3_AND8_NUM792_OUT));
      NOR2_X1 XNOR_5_3_AND8_NUM792 (.ZN (XNOR_5_3_AND8_NUM792_OUT), .A1 (XNOR_5_1_AND8_NUM792_OUT), .A2 (XNOR_5_2_AND8_NUM792_OUT));

      wire XNOR_6_1_AND8_NUM792_OUT, XNOR_6_2_AND8_NUM792_OUT, XNOR_6_3_AND8_NUM792_OUT;
      NOR2_X1 XNOR_6_1_AND8_NUM792 (.ZN (XNOR_6_1_AND8_NUM792_OUT), .A1 (XNOR_3_3_AND8_NUM792_OUT), .A2 (GND));
      NOR2_X1 XNOR_6_2_AND8_NUM792 (.ZN (XNOR_6_2_AND8_NUM792_OUT), .A1 (GND), .A2 (XNOR_4_3_AND8_NUM792_OUT));
      NOR2_X1 XNOR_6_3_AND8_NUM792 (.ZN (XNOR_6_3_AND8_NUM792_OUT), .A1 (XNOR_6_1_AND8_NUM792_OUT), .A2 (XNOR_6_2_AND8_NUM792_OUT));

      wire XNOR_7_1_AND8_NUM792_OUT, XNOR_7_2_AND8_NUM792_OUT;
      NOR2_X1 XNOR_7_1_AND8_NUM792 (.ZN (XNOR_7_1_AND8_NUM792_OUT), .A1 (XNOR_5_3_AND8_NUM792_OUT), .A2 (GND));
      NOR2_X1 XNOR_7_2_AND8_NUM792 (.ZN (XNOR_7_2_AND8_NUM792_OUT), .A1 (GND), .A2 (XNOR_6_3_AND8_NUM792_OUT));
      NOR2_X1 XNOR_7_3_AND8_NUM792 (.ZN (N2747), .A1 (XNOR_7_1_AND8_NUM792_OUT), .A2 (XNOR_7_2_AND8_NUM792_OUT));
      wire XNOR_1_1_AND8_NUM793_OUT, XNOR_1_2_AND8_NUM793_OUT, XNOR_1_3_AND8_NUM793_OUT;
      NOR2_X1 XNOR_1_1_AND8_NUM793 (.ZN (XNOR_1_1_AND8_NUM793_OUT), .A1 (N2606), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND8_NUM793 (.ZN (XNOR_1_2_AND8_NUM793_OUT), .A1 (GND), .A2 (N2549));
      NOR2_X1 XNOR_1_3_AND8_NUM793 (.ZN (XNOR_1_3_AND8_NUM793_OUT), .A1 (XNOR_1_1_AND8_NUM793_OUT), .A2 (XNOR_1_2_AND8_NUM793_OUT));

      wire XNOR_2_1_AND8_NUM793_OUT, XNOR_2_2_AND8_NUM793_OUT, XNOR_2_3_AND8_NUM793_OUT;
      NOR2_X1 XNOR_2_1_AND8_NUM793 (.ZN (XNOR_2_1_AND8_NUM793_OUT), .A1 (N2611), .A2 (GND));
      NOR2_X1 XNOR_2_2_AND8_NUM793 (.ZN (XNOR_2_2_AND8_NUM793_OUT), .A1 (GND), .A2 (N2614));
      NOR2_X1 XNOR_2_3_AND8_NUM793 (.ZN (XNOR_2_3_AND8_NUM793_OUT), .A1 (XNOR_2_1_AND8_NUM793_OUT), .A2 (XNOR_2_2_AND8_NUM793_OUT));

      wire XNOR_3_1_AND8_NUM793_OUT, XNOR_3_2_AND8_NUM793_OUT, XNOR_3_3_AND8_NUM793_OUT;
      NOR2_X1 XNOR_3_1_AND8_NUM793 (.ZN (XNOR_3_1_AND8_NUM793_OUT), .A1 (N2617), .A2 (GND));
      NOR2_X1 XNOR_3_2_AND8_NUM793 (.ZN (XNOR_3_2_AND8_NUM793_OUT), .A1 (GND), .A2 (N2620));
      NOR2_X1 XNOR_3_3_AND8_NUM793 (.ZN (XNOR_3_3_AND8_NUM793_OUT), .A1 (XNOR_3_1_AND8_NUM793_OUT), .A2 (XNOR_3_2_AND8_NUM793_OUT));

      wire XNOR_4_1_AND8_NUM793_OUT, XNOR_4_2_AND8_NUM793_OUT, XNOR_4_3_AND8_NUM793_OUT;
      NOR2_X1 XNOR_4_1_AND8_NUM793 (.ZN (XNOR_4_1_AND8_NUM793_OUT), .A1 (N2552), .A2 (GND));
      NOR2_X1 XNOR_4_2_AND8_NUM793 (.ZN (XNOR_4_2_AND8_NUM793_OUT), .A1 (GND), .A2 (N2555));
      NOR2_X1 XNOR_4_3_AND8_NUM793 (.ZN (XNOR_4_3_AND8_NUM793_OUT), .A1 (XNOR_4_1_AND8_NUM793_OUT), .A2 (XNOR_4_2_AND8_NUM793_OUT));

      wire XNOR_5_1_AND8_NUM793_OUT, XNOR_5_2_AND8_NUM793_OUT, XNOR_5_3_AND8_NUM793_OUT;
      NOR2_X1 XNOR_5_1_AND8_NUM793 (.ZN (XNOR_5_1_AND8_NUM793_OUT), .A1 (XNOR_1_3_AND8_NUM793_OUT), .A2 (GND));
      NOR2_X1 XNOR_5_2_AND8_NUM793 (.ZN (XNOR_5_2_AND8_NUM793_OUT), .A1 (GND), .A2 (XNOR_2_3_AND8_NUM793_OUT));
      NOR2_X1 XNOR_5_3_AND8_NUM793 (.ZN (XNOR_5_3_AND8_NUM793_OUT), .A1 (XNOR_5_1_AND8_NUM793_OUT), .A2 (XNOR_5_2_AND8_NUM793_OUT));

      wire XNOR_6_1_AND8_NUM793_OUT, XNOR_6_2_AND8_NUM793_OUT, XNOR_6_3_AND8_NUM793_OUT;
      NOR2_X1 XNOR_6_1_AND8_NUM793 (.ZN (XNOR_6_1_AND8_NUM793_OUT), .A1 (XNOR_3_3_AND8_NUM793_OUT), .A2 (GND));
      NOR2_X1 XNOR_6_2_AND8_NUM793 (.ZN (XNOR_6_2_AND8_NUM793_OUT), .A1 (GND), .A2 (XNOR_4_3_AND8_NUM793_OUT));
      NOR2_X1 XNOR_6_3_AND8_NUM793 (.ZN (XNOR_6_3_AND8_NUM793_OUT), .A1 (XNOR_6_1_AND8_NUM793_OUT), .A2 (XNOR_6_2_AND8_NUM793_OUT));

      wire XNOR_7_1_AND8_NUM793_OUT, XNOR_7_2_AND8_NUM793_OUT;
      NOR2_X1 XNOR_7_1_AND8_NUM793 (.ZN (XNOR_7_1_AND8_NUM793_OUT), .A1 (XNOR_5_3_AND8_NUM793_OUT), .A2 (GND));
      NOR2_X1 XNOR_7_2_AND8_NUM793 (.ZN (XNOR_7_2_AND8_NUM793_OUT), .A1 (GND), .A2 (XNOR_6_3_AND8_NUM793_OUT));
      NOR2_X1 XNOR_7_3_AND8_NUM793 (.ZN (N2750), .A1 (XNOR_7_1_AND8_NUM793_OUT), .A2 (XNOR_7_2_AND8_NUM793_OUT));
      wire XNOR_1_1_NAND2_NUM794_OUT, XNOR_1_2_NAND2_NUM794_OUT, XNOR_1_3_NAND2_NUM794_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM794 (.ZN (XNOR_1_1_NAND2_NUM794_OUT), .A1 (N2669), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM794 (.ZN (XNOR_1_2_NAND2_NUM794_OUT), .A1 (GND), .A2 (N2720));
      NOR2_X1 XNOR_1_3_NAND2_NUM794 (.ZN (XNOR_1_3_NAND2_NUM794_OUT), .A1 (XNOR_1_1_NAND2_NUM794_OUT), .A2 (XNOR_1_2_NAND2_NUM794_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM794 (.ZN (N2753), .A1 (XNOR_1_3_NAND2_NUM794_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM795_OUT, XNOR_1_2_NAND2_NUM795_OUT, XNOR_1_3_NAND2_NUM795_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM795 (.ZN (XNOR_1_1_NAND2_NUM795_OUT), .A1 (N2671), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM795 (.ZN (XNOR_1_2_NAND2_NUM795_OUT), .A1 (GND), .A2 (N2721));
      NOR2_X1 XNOR_1_3_NAND2_NUM795 (.ZN (XNOR_1_3_NAND2_NUM795_OUT), .A1 (XNOR_1_1_NAND2_NUM795_OUT), .A2 (XNOR_1_2_NAND2_NUM795_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM795 (.ZN (N2754), .A1 (XNOR_1_3_NAND2_NUM795_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM796_OUT, XNOR_1_2_NAND2_NUM796_OUT, XNOR_1_3_NAND2_NUM796_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM796 (.ZN (XNOR_1_1_NAND2_NUM796_OUT), .A1 (N2673), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM796 (.ZN (XNOR_1_2_NAND2_NUM796_OUT), .A1 (GND), .A2 (N2722));
      NOR2_X1 XNOR_1_3_NAND2_NUM796 (.ZN (XNOR_1_3_NAND2_NUM796_OUT), .A1 (XNOR_1_1_NAND2_NUM796_OUT), .A2 (XNOR_1_2_NAND2_NUM796_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM796 (.ZN (N2755), .A1 (XNOR_1_3_NAND2_NUM796_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM797_OUT, XNOR_1_2_NAND2_NUM797_OUT, XNOR_1_3_NAND2_NUM797_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM797 (.ZN (XNOR_1_1_NAND2_NUM797_OUT), .A1 (N2675), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM797 (.ZN (XNOR_1_2_NAND2_NUM797_OUT), .A1 (GND), .A2 (N2723));
      NOR2_X1 XNOR_1_3_NAND2_NUM797 (.ZN (XNOR_1_3_NAND2_NUM797_OUT), .A1 (XNOR_1_1_NAND2_NUM797_OUT), .A2 (XNOR_1_2_NAND2_NUM797_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM797 (.ZN (N2756), .A1 (XNOR_1_3_NAND2_NUM797_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM798_OUT, XNOR_1_2_NAND2_NUM798_OUT, XNOR_1_3_NAND2_NUM798_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM798 (.ZN (XNOR_1_1_NAND2_NUM798_OUT), .A1 (N355), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM798 (.ZN (XNOR_1_2_NAND2_NUM798_OUT), .A1 (GND), .A2 (N2725));
      NOR2_X1 XNOR_1_3_NAND2_NUM798 (.ZN (XNOR_1_3_NAND2_NUM798_OUT), .A1 (XNOR_1_1_NAND2_NUM798_OUT), .A2 (XNOR_1_2_NAND2_NUM798_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM798 (.ZN (N2757), .A1 (XNOR_1_3_NAND2_NUM798_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM799_OUT, XNOR_1_2_NAND2_NUM799_OUT, XNOR_1_3_NAND2_NUM799_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM799 (.ZN (XNOR_1_1_NAND2_NUM799_OUT), .A1 (N358), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM799 (.ZN (XNOR_1_2_NAND2_NUM799_OUT), .A1 (GND), .A2 (N2727));
      NOR2_X1 XNOR_1_3_NAND2_NUM799 (.ZN (XNOR_1_3_NAND2_NUM799_OUT), .A1 (XNOR_1_1_NAND2_NUM799_OUT), .A2 (XNOR_1_2_NAND2_NUM799_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM799 (.ZN (N2758), .A1 (XNOR_1_3_NAND2_NUM799_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM800_OUT, XNOR_1_2_NAND2_NUM800_OUT, XNOR_1_3_NAND2_NUM800_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM800 (.ZN (XNOR_1_1_NAND2_NUM800_OUT), .A1 (N361), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM800 (.ZN (XNOR_1_2_NAND2_NUM800_OUT), .A1 (GND), .A2 (N2729));
      NOR2_X1 XNOR_1_3_NAND2_NUM800 (.ZN (XNOR_1_3_NAND2_NUM800_OUT), .A1 (XNOR_1_1_NAND2_NUM800_OUT), .A2 (XNOR_1_2_NAND2_NUM800_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM800 (.ZN (N2759), .A1 (XNOR_1_3_NAND2_NUM800_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM801_OUT, XNOR_1_2_NAND2_NUM801_OUT, XNOR_1_3_NAND2_NUM801_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM801 (.ZN (XNOR_1_1_NAND2_NUM801_OUT), .A1 (N364), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM801 (.ZN (XNOR_1_2_NAND2_NUM801_OUT), .A1 (GND), .A2 (N2731));
      NOR2_X1 XNOR_1_3_NAND2_NUM801 (.ZN (XNOR_1_3_NAND2_NUM801_OUT), .A1 (XNOR_1_1_NAND2_NUM801_OUT), .A2 (XNOR_1_2_NAND2_NUM801_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM801 (.ZN (N2760), .A1 (XNOR_1_3_NAND2_NUM801_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM802_OUT, XNOR_1_2_NAND2_NUM802_OUT, XNOR_1_3_NAND2_NUM802_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM802 (.ZN (XNOR_1_1_NAND2_NUM802_OUT), .A1 (N367), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM802 (.ZN (XNOR_1_2_NAND2_NUM802_OUT), .A1 (GND), .A2 (N2733));
      NOR2_X1 XNOR_1_3_NAND2_NUM802 (.ZN (XNOR_1_3_NAND2_NUM802_OUT), .A1 (XNOR_1_1_NAND2_NUM802_OUT), .A2 (XNOR_1_2_NAND2_NUM802_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM802 (.ZN (N2761), .A1 (XNOR_1_3_NAND2_NUM802_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM803_OUT, XNOR_1_2_NAND2_NUM803_OUT, XNOR_1_3_NAND2_NUM803_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM803 (.ZN (XNOR_1_1_NAND2_NUM803_OUT), .A1 (N2682), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM803 (.ZN (XNOR_1_2_NAND2_NUM803_OUT), .A1 (GND), .A2 (N2734));
      NOR2_X1 XNOR_1_3_NAND2_NUM803 (.ZN (XNOR_1_3_NAND2_NUM803_OUT), .A1 (XNOR_1_1_NAND2_NUM803_OUT), .A2 (XNOR_1_2_NAND2_NUM803_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM803 (.ZN (N2762), .A1 (XNOR_1_3_NAND2_NUM803_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM804_OUT, XNOR_1_2_NAND2_NUM804_OUT, XNOR_1_3_NAND2_NUM804_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM804 (.ZN (XNOR_1_1_NAND2_NUM804_OUT), .A1 (N373), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM804 (.ZN (XNOR_1_2_NAND2_NUM804_OUT), .A1 (GND), .A2 (N2736));
      NOR2_X1 XNOR_1_3_NAND2_NUM804 (.ZN (XNOR_1_3_NAND2_NUM804_OUT), .A1 (XNOR_1_1_NAND2_NUM804_OUT), .A2 (XNOR_1_2_NAND2_NUM804_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM804 (.ZN (N2763), .A1 (XNOR_1_3_NAND2_NUM804_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM805_OUT, XNOR_1_2_NAND2_NUM805_OUT, XNOR_1_3_NAND2_NUM805_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM805 (.ZN (XNOR_1_1_NAND2_NUM805_OUT), .A1 (N376), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM805 (.ZN (XNOR_1_2_NAND2_NUM805_OUT), .A1 (GND), .A2 (N2738));
      NOR2_X1 XNOR_1_3_NAND2_NUM805 (.ZN (XNOR_1_3_NAND2_NUM805_OUT), .A1 (XNOR_1_1_NAND2_NUM805_OUT), .A2 (XNOR_1_2_NAND2_NUM805_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM805 (.ZN (N2764), .A1 (XNOR_1_3_NAND2_NUM805_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM806_OUT, XNOR_1_2_NAND2_NUM806_OUT, XNOR_1_3_NAND2_NUM806_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM806 (.ZN (XNOR_1_1_NAND2_NUM806_OUT), .A1 (N379), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM806 (.ZN (XNOR_1_2_NAND2_NUM806_OUT), .A1 (GND), .A2 (N2740));
      NOR2_X1 XNOR_1_3_NAND2_NUM806 (.ZN (XNOR_1_3_NAND2_NUM806_OUT), .A1 (XNOR_1_1_NAND2_NUM806_OUT), .A2 (XNOR_1_2_NAND2_NUM806_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM806 (.ZN (N2765), .A1 (XNOR_1_3_NAND2_NUM806_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM807_OUT, XNOR_1_2_NAND2_NUM807_OUT, XNOR_1_3_NAND2_NUM807_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM807 (.ZN (XNOR_1_1_NAND2_NUM807_OUT), .A1 (N382), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM807 (.ZN (XNOR_1_2_NAND2_NUM807_OUT), .A1 (GND), .A2 (N2742));
      NOR2_X1 XNOR_1_3_NAND2_NUM807 (.ZN (XNOR_1_3_NAND2_NUM807_OUT), .A1 (XNOR_1_1_NAND2_NUM807_OUT), .A2 (XNOR_1_2_NAND2_NUM807_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM807 (.ZN (N2766), .A1 (XNOR_1_3_NAND2_NUM807_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM808_OUT, XNOR_1_2_NAND2_NUM808_OUT, XNOR_1_3_NAND2_NUM808_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM808 (.ZN (XNOR_1_1_NAND2_NUM808_OUT), .A1 (N2688), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM808 (.ZN (XNOR_1_2_NAND2_NUM808_OUT), .A1 (GND), .A2 (N2743));
      NOR2_X1 XNOR_1_3_NAND2_NUM808 (.ZN (XNOR_1_3_NAND2_NUM808_OUT), .A1 (XNOR_1_1_NAND2_NUM808_OUT), .A2 (XNOR_1_2_NAND2_NUM808_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM808 (.ZN (N2767), .A1 (XNOR_1_3_NAND2_NUM808_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM809_OUT, XNOR_1_2_NAND2_NUM809_OUT, XNOR_1_3_NAND2_NUM809_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM809 (.ZN (XNOR_1_1_NAND2_NUM809_OUT), .A1 (N2690), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM809 (.ZN (XNOR_1_2_NAND2_NUM809_OUT), .A1 (GND), .A2 (N2744));
      NOR2_X1 XNOR_1_3_NAND2_NUM809 (.ZN (XNOR_1_3_NAND2_NUM809_OUT), .A1 (XNOR_1_1_NAND2_NUM809_OUT), .A2 (XNOR_1_2_NAND2_NUM809_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM809 (.ZN (N2768), .A1 (XNOR_1_3_NAND2_NUM809_OUT), .A2 (GND));
      wire XNOR_1_1_AND2_NUM810_OUT, XNOR_1_2_AND2_NUM810_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM810 (.ZN (XNOR_1_1_AND2_NUM810_OUT), .A1 (N2745), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM810 (.ZN (XNOR_1_2_AND2_NUM810_OUT), .A1 (GND), .A2 (N275));
      NOR2_X1 XNOR_1_3_AND2_NUM810 (.ZN (N2773), .A1 (XNOR_1_1_AND2_NUM810_OUT), .A2 (XNOR_1_2_AND2_NUM810_OUT));
      wire XNOR_1_1_AND2_NUM811_OUT, XNOR_1_2_AND2_NUM811_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM811 (.ZN (XNOR_1_1_AND2_NUM811_OUT), .A1 (N2746), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM811 (.ZN (XNOR_1_2_AND2_NUM811_OUT), .A1 (GND), .A2 (N276));
      NOR2_X1 XNOR_1_3_AND2_NUM811 (.ZN (N2776), .A1 (XNOR_1_1_AND2_NUM811_OUT), .A2 (XNOR_1_2_AND2_NUM811_OUT));
      wire XNOR_1_1_NAND2_NUM812_OUT, XNOR_1_2_NAND2_NUM812_OUT, XNOR_1_3_NAND2_NUM812_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM812 (.ZN (XNOR_1_1_NAND2_NUM812_OUT), .A1 (N2724), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM812 (.ZN (XNOR_1_2_NAND2_NUM812_OUT), .A1 (GND), .A2 (N2757));
      NOR2_X1 XNOR_1_3_NAND2_NUM812 (.ZN (XNOR_1_3_NAND2_NUM812_OUT), .A1 (XNOR_1_1_NAND2_NUM812_OUT), .A2 (XNOR_1_2_NAND2_NUM812_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM812 (.ZN (N2779), .A1 (XNOR_1_3_NAND2_NUM812_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM813_OUT, XNOR_1_2_NAND2_NUM813_OUT, XNOR_1_3_NAND2_NUM813_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM813 (.ZN (XNOR_1_1_NAND2_NUM813_OUT), .A1 (N2726), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM813 (.ZN (XNOR_1_2_NAND2_NUM813_OUT), .A1 (GND), .A2 (N2758));
      NOR2_X1 XNOR_1_3_NAND2_NUM813 (.ZN (XNOR_1_3_NAND2_NUM813_OUT), .A1 (XNOR_1_1_NAND2_NUM813_OUT), .A2 (XNOR_1_2_NAND2_NUM813_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM813 (.ZN (N2780), .A1 (XNOR_1_3_NAND2_NUM813_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM814_OUT, XNOR_1_2_NAND2_NUM814_OUT, XNOR_1_3_NAND2_NUM814_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM814 (.ZN (XNOR_1_1_NAND2_NUM814_OUT), .A1 (N2728), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM814 (.ZN (XNOR_1_2_NAND2_NUM814_OUT), .A1 (GND), .A2 (N2759));
      NOR2_X1 XNOR_1_3_NAND2_NUM814 (.ZN (XNOR_1_3_NAND2_NUM814_OUT), .A1 (XNOR_1_1_NAND2_NUM814_OUT), .A2 (XNOR_1_2_NAND2_NUM814_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM814 (.ZN (N2781), .A1 (XNOR_1_3_NAND2_NUM814_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM815_OUT, XNOR_1_2_NAND2_NUM815_OUT, XNOR_1_3_NAND2_NUM815_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM815 (.ZN (XNOR_1_1_NAND2_NUM815_OUT), .A1 (N2730), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM815 (.ZN (XNOR_1_2_NAND2_NUM815_OUT), .A1 (GND), .A2 (N2760));
      NOR2_X1 XNOR_1_3_NAND2_NUM815 (.ZN (XNOR_1_3_NAND2_NUM815_OUT), .A1 (XNOR_1_1_NAND2_NUM815_OUT), .A2 (XNOR_1_2_NAND2_NUM815_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM815 (.ZN (N2782), .A1 (XNOR_1_3_NAND2_NUM815_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM816_OUT, XNOR_1_2_NAND2_NUM816_OUT, XNOR_1_3_NAND2_NUM816_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM816 (.ZN (XNOR_1_1_NAND2_NUM816_OUT), .A1 (N2732), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM816 (.ZN (XNOR_1_2_NAND2_NUM816_OUT), .A1 (GND), .A2 (N2761));
      NOR2_X1 XNOR_1_3_NAND2_NUM816 (.ZN (XNOR_1_3_NAND2_NUM816_OUT), .A1 (XNOR_1_1_NAND2_NUM816_OUT), .A2 (XNOR_1_2_NAND2_NUM816_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM816 (.ZN (N2783), .A1 (XNOR_1_3_NAND2_NUM816_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM817_OUT, XNOR_1_2_NAND2_NUM817_OUT, XNOR_1_3_NAND2_NUM817_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM817 (.ZN (XNOR_1_1_NAND2_NUM817_OUT), .A1 (N2735), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM817 (.ZN (XNOR_1_2_NAND2_NUM817_OUT), .A1 (GND), .A2 (N2763));
      NOR2_X1 XNOR_1_3_NAND2_NUM817 (.ZN (XNOR_1_3_NAND2_NUM817_OUT), .A1 (XNOR_1_1_NAND2_NUM817_OUT), .A2 (XNOR_1_2_NAND2_NUM817_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM817 (.ZN (N2784), .A1 (XNOR_1_3_NAND2_NUM817_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM818_OUT, XNOR_1_2_NAND2_NUM818_OUT, XNOR_1_3_NAND2_NUM818_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM818 (.ZN (XNOR_1_1_NAND2_NUM818_OUT), .A1 (N2737), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM818 (.ZN (XNOR_1_2_NAND2_NUM818_OUT), .A1 (GND), .A2 (N2764));
      NOR2_X1 XNOR_1_3_NAND2_NUM818 (.ZN (XNOR_1_3_NAND2_NUM818_OUT), .A1 (XNOR_1_1_NAND2_NUM818_OUT), .A2 (XNOR_1_2_NAND2_NUM818_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM818 (.ZN (N2785), .A1 (XNOR_1_3_NAND2_NUM818_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM819_OUT, XNOR_1_2_NAND2_NUM819_OUT, XNOR_1_3_NAND2_NUM819_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM819 (.ZN (XNOR_1_1_NAND2_NUM819_OUT), .A1 (N2739), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM819 (.ZN (XNOR_1_2_NAND2_NUM819_OUT), .A1 (GND), .A2 (N2765));
      NOR2_X1 XNOR_1_3_NAND2_NUM819 (.ZN (XNOR_1_3_NAND2_NUM819_OUT), .A1 (XNOR_1_1_NAND2_NUM819_OUT), .A2 (XNOR_1_2_NAND2_NUM819_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM819 (.ZN (N2786), .A1 (XNOR_1_3_NAND2_NUM819_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM820_OUT, XNOR_1_2_NAND2_NUM820_OUT, XNOR_1_3_NAND2_NUM820_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM820 (.ZN (XNOR_1_1_NAND2_NUM820_OUT), .A1 (N2741), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM820 (.ZN (XNOR_1_2_NAND2_NUM820_OUT), .A1 (GND), .A2 (N2766));
      NOR2_X1 XNOR_1_3_NAND2_NUM820 (.ZN (XNOR_1_3_NAND2_NUM820_OUT), .A1 (XNOR_1_1_NAND2_NUM820_OUT), .A2 (XNOR_1_2_NAND2_NUM820_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM820 (.ZN (N2787), .A1 (XNOR_1_3_NAND2_NUM820_OUT), .A2 (GND));
      wire XNOR_1_1_AND3_NUM821_OUT, XNOR_1_2_AND3_NUM821_OUT, XNOR_1_3_AND3_NUM821_OUT;
      NOR2_X1 XNOR_1_1_AND3_NUM821 (.ZN (XNOR_1_1_AND3_NUM821_OUT), .A1 (N2747), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND3_NUM821 (.ZN (XNOR_1_2_AND3_NUM821_OUT), .A1 (GND), .A2 (N2750));
      NOR2_X1 XNOR_1_3_AND3_NUM821 (.ZN (XNOR_1_3_AND3_NUM821_OUT), .A1 (XNOR_1_1_AND3_NUM821_OUT), .A2 (XNOR_1_2_AND3_NUM821_OUT));

      wire XNOR_2_1_AND3_NUM821_OUT, XNOR_2_2_AND3_NUM821_OUT;
      NOR2_X1 XNOR_2_1_AND3_NUM821 (.ZN (XNOR_2_1_AND3_NUM821_OUT), .A1 (N2710), .A2 (GND));
      NOR2_X1 XNOR_2_2_AND3_NUM821 (.ZN (XNOR_2_2_AND3_NUM821_OUT), .A1 (GND), .A2 (XNOR_1_3_AND3_NUM821_OUT));
      NOR2_X1 XNOR_2_3_AND3_NUM821 (.ZN (N2788), .A1 (XNOR_2_1_AND3_NUM821_OUT), .A2 (XNOR_2_2_AND3_NUM821_OUT));
      wire XNOR_1_1_NAND2_NUM822_OUT, XNOR_1_2_NAND2_NUM822_OUT, XNOR_1_3_NAND2_NUM822_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM822 (.ZN (XNOR_1_1_NAND2_NUM822_OUT), .A1 (N2747), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM822 (.ZN (XNOR_1_2_NAND2_NUM822_OUT), .A1 (GND), .A2 (N2750));
      NOR2_X1 XNOR_1_3_NAND2_NUM822 (.ZN (XNOR_1_3_NAND2_NUM822_OUT), .A1 (XNOR_1_1_NAND2_NUM822_OUT), .A2 (XNOR_1_2_NAND2_NUM822_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM822 (.ZN (N2789), .A1 (XNOR_1_3_NAND2_NUM822_OUT), .A2 (GND));
      wire XNOR_1_1_AND4_NUM823_OUT, XNOR_1_2_AND4_NUM823_OUT, XNOR_1_3_AND4_NUM823_OUT;
      NOR2_X1 XNOR_1_1_AND4_NUM823 (.ZN (XNOR_1_1_AND4_NUM823_OUT), .A1 (N338), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND4_NUM823 (.ZN (XNOR_1_2_AND4_NUM823_OUT), .A1 (GND), .A2 (N2279));
      NOR2_X1 XNOR_1_3_AND4_NUM823 (.ZN (XNOR_1_3_AND4_NUM823_OUT), .A1 (XNOR_1_1_AND4_NUM823_OUT), .A2 (XNOR_1_2_AND4_NUM823_OUT));

      wire XNOR_2_1_AND4_NUM823_OUT, XNOR_2_2_AND4_NUM823_OUT, XNOR_2_3_AND4_NUM823_OUT;
      NOR2_X1 XNOR_2_1_AND4_NUM823 (.ZN (XNOR_2_1_AND4_NUM823_OUT), .A1 (N99), .A2 (GND));
      NOR2_X1 XNOR_2_2_AND4_NUM823 (.ZN (XNOR_2_2_AND4_NUM823_OUT), .A1 (GND), .A2 (N2788));
      NOR2_X1 XNOR_2_3_AND4_NUM823 (.ZN (XNOR_2_3_AND4_NUM823_OUT), .A1 (XNOR_2_1_AND4_NUM823_OUT), .A2 (XNOR_2_2_AND4_NUM823_OUT));

      wire XNOR_3_1_AND4_NUM823_OUT, XNOR_3_2_AND4_NUM823_OUT;
      NOR2_X1 XNOR_3_1_AND4_NUM823 (.ZN (XNOR_3_1_AND4_NUM823_OUT), .A1 (XNOR_1_3_AND4_NUM823_OUT), .A2 (GND));
      NOR2_X1 XNOR_3_2_AND4_NUM823 (.ZN (XNOR_3_2_AND4_NUM823_OUT), .A1 (GND), .A2 (XNOR_2_3_AND4_NUM823_OUT));
      NOR2_X1 XNOR_3_3_AND4_NUM823 (.ZN (N2800), .A1 (XNOR_3_1_AND4_NUM823_OUT), .A2 (XNOR_3_2_AND4_NUM823_OUT));
      wire XNOR_1_1_NAND2_NUM824_OUT, XNOR_1_2_NAND2_NUM824_OUT, XNOR_1_3_NAND2_NUM824_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM824 (.ZN (XNOR_1_1_NAND2_NUM824_OUT), .A1 (N2773), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM824 (.ZN (XNOR_1_2_NAND2_NUM824_OUT), .A1 (GND), .A2 (N2018));
      NOR2_X1 XNOR_1_3_NAND2_NUM824 (.ZN (XNOR_1_3_NAND2_NUM824_OUT), .A1 (XNOR_1_1_NAND2_NUM824_OUT), .A2 (XNOR_1_2_NAND2_NUM824_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM824 (.ZN (N2807), .A1 (XNOR_1_3_NAND2_NUM824_OUT), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM825 (.ZN (N2808), .A1 (N2773), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM826_OUT, XNOR_1_2_NAND2_NUM826_OUT, XNOR_1_3_NAND2_NUM826_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM826 (.ZN (XNOR_1_1_NAND2_NUM826_OUT), .A1 (N2776), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM826 (.ZN (XNOR_1_2_NAND2_NUM826_OUT), .A1 (GND), .A2 (N2019));
      NOR2_X1 XNOR_1_3_NAND2_NUM826 (.ZN (XNOR_1_3_NAND2_NUM826_OUT), .A1 (XNOR_1_1_NAND2_NUM826_OUT), .A2 (XNOR_1_2_NAND2_NUM826_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM826 (.ZN (N2809), .A1 (XNOR_1_3_NAND2_NUM826_OUT), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM827 (.ZN (N2810), .A1 (N2776), .A2 (GND));
      NOR2_X1 XNOR_NOR2_NUM828 (.ZN (N2811), .A1 (N2384), .A2 (N2800));
      wire XNOR_1_1_AND3_NUM829_OUT, XNOR_1_2_AND3_NUM829_OUT, XNOR_1_3_AND3_NUM829_OUT;
      NOR2_X1 XNOR_1_1_AND3_NUM829 (.ZN (XNOR_1_1_AND3_NUM829_OUT), .A1 (N897), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND3_NUM829 (.ZN (XNOR_1_2_AND3_NUM829_OUT), .A1 (GND), .A2 (N283));
      NOR2_X1 XNOR_1_3_AND3_NUM829 (.ZN (XNOR_1_3_AND3_NUM829_OUT), .A1 (XNOR_1_1_AND3_NUM829_OUT), .A2 (XNOR_1_2_AND3_NUM829_OUT));

      wire XNOR_2_1_AND3_NUM829_OUT, XNOR_2_2_AND3_NUM829_OUT;
      NOR2_X1 XNOR_2_1_AND3_NUM829 (.ZN (XNOR_2_1_AND3_NUM829_OUT), .A1 (N2789), .A2 (GND));
      NOR2_X1 XNOR_2_2_AND3_NUM829 (.ZN (XNOR_2_2_AND3_NUM829_OUT), .A1 (GND), .A2 (XNOR_1_3_AND3_NUM829_OUT));
      NOR2_X1 XNOR_2_3_AND3_NUM829 (.ZN (N2812), .A1 (XNOR_2_1_AND3_NUM829_OUT), .A2 (XNOR_2_2_AND3_NUM829_OUT));
      wire XNOR_1_1_AND3_NUM830_OUT, XNOR_1_2_AND3_NUM830_OUT, XNOR_1_3_AND3_NUM830_OUT;
      NOR2_X1 XNOR_1_1_AND3_NUM830 (.ZN (XNOR_1_1_AND3_NUM830_OUT), .A1 (N76), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND3_NUM830 (.ZN (XNOR_1_2_AND3_NUM830_OUT), .A1 (GND), .A2 (N283));
      NOR2_X1 XNOR_1_3_AND3_NUM830 (.ZN (XNOR_1_3_AND3_NUM830_OUT), .A1 (XNOR_1_1_AND3_NUM830_OUT), .A2 (XNOR_1_2_AND3_NUM830_OUT));

      wire XNOR_2_1_AND3_NUM830_OUT, XNOR_2_2_AND3_NUM830_OUT;
      NOR2_X1 XNOR_2_1_AND3_NUM830 (.ZN (XNOR_2_1_AND3_NUM830_OUT), .A1 (N2789), .A2 (GND));
      NOR2_X1 XNOR_2_2_AND3_NUM830 (.ZN (XNOR_2_2_AND3_NUM830_OUT), .A1 (GND), .A2 (XNOR_1_3_AND3_NUM830_OUT));
      NOR2_X1 XNOR_2_3_AND3_NUM830 (.ZN (N2815), .A1 (XNOR_2_1_AND3_NUM830_OUT), .A2 (XNOR_2_2_AND3_NUM830_OUT));
      wire XNOR_1_1_AND3_NUM831_OUT, XNOR_1_2_AND3_NUM831_OUT, XNOR_1_3_AND3_NUM831_OUT;
      NOR2_X1 XNOR_1_1_AND3_NUM831 (.ZN (XNOR_1_1_AND3_NUM831_OUT), .A1 (N82), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND3_NUM831 (.ZN (XNOR_1_2_AND3_NUM831_OUT), .A1 (GND), .A2 (N283));
      NOR2_X1 XNOR_1_3_AND3_NUM831 (.ZN (XNOR_1_3_AND3_NUM831_OUT), .A1 (XNOR_1_1_AND3_NUM831_OUT), .A2 (XNOR_1_2_AND3_NUM831_OUT));

      wire XNOR_2_1_AND3_NUM831_OUT, XNOR_2_2_AND3_NUM831_OUT;
      NOR2_X1 XNOR_2_1_AND3_NUM831 (.ZN (XNOR_2_1_AND3_NUM831_OUT), .A1 (N2789), .A2 (GND));
      NOR2_X1 XNOR_2_2_AND3_NUM831 (.ZN (XNOR_2_2_AND3_NUM831_OUT), .A1 (GND), .A2 (XNOR_1_3_AND3_NUM831_OUT));
      NOR2_X1 XNOR_2_3_AND3_NUM831 (.ZN (N2818), .A1 (XNOR_2_1_AND3_NUM831_OUT), .A2 (XNOR_2_2_AND3_NUM831_OUT));
      wire XNOR_1_1_AND3_NUM832_OUT, XNOR_1_2_AND3_NUM832_OUT, XNOR_1_3_AND3_NUM832_OUT;
      NOR2_X1 XNOR_1_1_AND3_NUM832 (.ZN (XNOR_1_1_AND3_NUM832_OUT), .A1 (N85), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND3_NUM832 (.ZN (XNOR_1_2_AND3_NUM832_OUT), .A1 (GND), .A2 (N283));
      NOR2_X1 XNOR_1_3_AND3_NUM832 (.ZN (XNOR_1_3_AND3_NUM832_OUT), .A1 (XNOR_1_1_AND3_NUM832_OUT), .A2 (XNOR_1_2_AND3_NUM832_OUT));

      wire XNOR_2_1_AND3_NUM832_OUT, XNOR_2_2_AND3_NUM832_OUT;
      NOR2_X1 XNOR_2_1_AND3_NUM832 (.ZN (XNOR_2_1_AND3_NUM832_OUT), .A1 (N2789), .A2 (GND));
      NOR2_X1 XNOR_2_2_AND3_NUM832 (.ZN (XNOR_2_2_AND3_NUM832_OUT), .A1 (GND), .A2 (XNOR_1_3_AND3_NUM832_OUT));
      NOR2_X1 XNOR_2_3_AND3_NUM832 (.ZN (N2821), .A1 (XNOR_2_1_AND3_NUM832_OUT), .A2 (XNOR_2_2_AND3_NUM832_OUT));
      wire XNOR_1_1_AND3_NUM833_OUT, XNOR_1_2_AND3_NUM833_OUT, XNOR_1_3_AND3_NUM833_OUT;
      NOR2_X1 XNOR_1_1_AND3_NUM833 (.ZN (XNOR_1_1_AND3_NUM833_OUT), .A1 (N898), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND3_NUM833 (.ZN (XNOR_1_2_AND3_NUM833_OUT), .A1 (GND), .A2 (N283));
      NOR2_X1 XNOR_1_3_AND3_NUM833 (.ZN (XNOR_1_3_AND3_NUM833_OUT), .A1 (XNOR_1_1_AND3_NUM833_OUT), .A2 (XNOR_1_2_AND3_NUM833_OUT));

      wire XNOR_2_1_AND3_NUM833_OUT, XNOR_2_2_AND3_NUM833_OUT;
      NOR2_X1 XNOR_2_1_AND3_NUM833 (.ZN (XNOR_2_1_AND3_NUM833_OUT), .A1 (N2789), .A2 (GND));
      NOR2_X1 XNOR_2_2_AND3_NUM833 (.ZN (XNOR_2_2_AND3_NUM833_OUT), .A1 (GND), .A2 (XNOR_1_3_AND3_NUM833_OUT));
      NOR2_X1 XNOR_2_3_AND3_NUM833 (.ZN (N2824), .A1 (XNOR_2_1_AND3_NUM833_OUT), .A2 (XNOR_2_2_AND3_NUM833_OUT));
      wire XNOR_1_1_NAND2_NUM834_OUT, XNOR_1_2_NAND2_NUM834_OUT, XNOR_1_3_NAND2_NUM834_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM834 (.ZN (XNOR_1_1_NAND2_NUM834_OUT), .A1 (N1965), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM834 (.ZN (XNOR_1_2_NAND2_NUM834_OUT), .A1 (GND), .A2 (N2808));
      NOR2_X1 XNOR_1_3_NAND2_NUM834 (.ZN (XNOR_1_3_NAND2_NUM834_OUT), .A1 (XNOR_1_1_NAND2_NUM834_OUT), .A2 (XNOR_1_2_NAND2_NUM834_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM834 (.ZN (N2827), .A1 (XNOR_1_3_NAND2_NUM834_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM835_OUT, XNOR_1_2_NAND2_NUM835_OUT, XNOR_1_3_NAND2_NUM835_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM835 (.ZN (XNOR_1_1_NAND2_NUM835_OUT), .A1 (N1968), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM835 (.ZN (XNOR_1_2_NAND2_NUM835_OUT), .A1 (GND), .A2 (N2810));
      NOR2_X1 XNOR_1_3_NAND2_NUM835 (.ZN (XNOR_1_3_NAND2_NUM835_OUT), .A1 (XNOR_1_1_NAND2_NUM835_OUT), .A2 (XNOR_1_2_NAND2_NUM835_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM835 (.ZN (N2828), .A1 (XNOR_1_3_NAND2_NUM835_OUT), .A2 (GND));
      wire XNOR_1_1_AND3_NUM836_OUT, XNOR_1_2_AND3_NUM836_OUT, XNOR_1_3_AND3_NUM836_OUT;
      NOR2_X1 XNOR_1_1_AND3_NUM836 (.ZN (XNOR_1_1_AND3_NUM836_OUT), .A1 (N79), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND3_NUM836 (.ZN (XNOR_1_2_AND3_NUM836_OUT), .A1 (GND), .A2 (N283));
      NOR2_X1 XNOR_1_3_AND3_NUM836 (.ZN (XNOR_1_3_AND3_NUM836_OUT), .A1 (XNOR_1_1_AND3_NUM836_OUT), .A2 (XNOR_1_2_AND3_NUM836_OUT));

      wire XNOR_2_1_AND3_NUM836_OUT, XNOR_2_2_AND3_NUM836_OUT;
      NOR2_X1 XNOR_2_1_AND3_NUM836 (.ZN (XNOR_2_1_AND3_NUM836_OUT), .A1 (N2789), .A2 (GND));
      NOR2_X1 XNOR_2_2_AND3_NUM836 (.ZN (XNOR_2_2_AND3_NUM836_OUT), .A1 (GND), .A2 (XNOR_1_3_AND3_NUM836_OUT));
      NOR2_X1 XNOR_2_3_AND3_NUM836 (.ZN (N2829), .A1 (XNOR_2_1_AND3_NUM836_OUT), .A2 (XNOR_2_2_AND3_NUM836_OUT));
      wire XNOR_1_1_NAND2_NUM837_OUT, XNOR_1_2_NAND2_NUM837_OUT, XNOR_1_3_NAND2_NUM837_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM837 (.ZN (XNOR_1_1_NAND2_NUM837_OUT), .A1 (N2807), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM837 (.ZN (XNOR_1_2_NAND2_NUM837_OUT), .A1 (GND), .A2 (N2827));
      NOR2_X1 XNOR_1_3_NAND2_NUM837 (.ZN (XNOR_1_3_NAND2_NUM837_OUT), .A1 (XNOR_1_1_NAND2_NUM837_OUT), .A2 (XNOR_1_2_NAND2_NUM837_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM837 (.ZN (N2843), .A1 (XNOR_1_3_NAND2_NUM837_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM838_OUT, XNOR_1_2_NAND2_NUM838_OUT, XNOR_1_3_NAND2_NUM838_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM838 (.ZN (XNOR_1_1_NAND2_NUM838_OUT), .A1 (N2809), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM838 (.ZN (XNOR_1_2_NAND2_NUM838_OUT), .A1 (GND), .A2 (N2828));
      NOR2_X1 XNOR_1_3_NAND2_NUM838 (.ZN (XNOR_1_3_NAND2_NUM838_OUT), .A1 (XNOR_1_1_NAND2_NUM838_OUT), .A2 (XNOR_1_2_NAND2_NUM838_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM838 (.ZN (N2846), .A1 (XNOR_1_3_NAND2_NUM838_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM839_OUT, XNOR_1_2_NAND2_NUM839_OUT, XNOR_1_3_NAND2_NUM839_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM839 (.ZN (XNOR_1_1_NAND2_NUM839_OUT), .A1 (N2812), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM839 (.ZN (XNOR_1_2_NAND2_NUM839_OUT), .A1 (GND), .A2 (N2076));
      NOR2_X1 XNOR_1_3_NAND2_NUM839 (.ZN (XNOR_1_3_NAND2_NUM839_OUT), .A1 (XNOR_1_1_NAND2_NUM839_OUT), .A2 (XNOR_1_2_NAND2_NUM839_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM839 (.ZN (N2850), .A1 (XNOR_1_3_NAND2_NUM839_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM840_OUT, XNOR_1_2_NAND2_NUM840_OUT, XNOR_1_3_NAND2_NUM840_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM840 (.ZN (XNOR_1_1_NAND2_NUM840_OUT), .A1 (N2815), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM840 (.ZN (XNOR_1_2_NAND2_NUM840_OUT), .A1 (GND), .A2 (N2077));
      NOR2_X1 XNOR_1_3_NAND2_NUM840 (.ZN (XNOR_1_3_NAND2_NUM840_OUT), .A1 (XNOR_1_1_NAND2_NUM840_OUT), .A2 (XNOR_1_2_NAND2_NUM840_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM840 (.ZN (N2851), .A1 (XNOR_1_3_NAND2_NUM840_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM841_OUT, XNOR_1_2_NAND2_NUM841_OUT, XNOR_1_3_NAND2_NUM841_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM841 (.ZN (XNOR_1_1_NAND2_NUM841_OUT), .A1 (N2818), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM841 (.ZN (XNOR_1_2_NAND2_NUM841_OUT), .A1 (GND), .A2 (N1915));
      NOR2_X1 XNOR_1_3_NAND2_NUM841 (.ZN (XNOR_1_3_NAND2_NUM841_OUT), .A1 (XNOR_1_1_NAND2_NUM841_OUT), .A2 (XNOR_1_2_NAND2_NUM841_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM841 (.ZN (N2852), .A1 (XNOR_1_3_NAND2_NUM841_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM842_OUT, XNOR_1_2_NAND2_NUM842_OUT, XNOR_1_3_NAND2_NUM842_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM842 (.ZN (XNOR_1_1_NAND2_NUM842_OUT), .A1 (N2821), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM842 (.ZN (XNOR_1_2_NAND2_NUM842_OUT), .A1 (GND), .A2 (N1857));
      NOR2_X1 XNOR_1_3_NAND2_NUM842 (.ZN (XNOR_1_3_NAND2_NUM842_OUT), .A1 (XNOR_1_1_NAND2_NUM842_OUT), .A2 (XNOR_1_2_NAND2_NUM842_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM842 (.ZN (N2853), .A1 (XNOR_1_3_NAND2_NUM842_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM843_OUT, XNOR_1_2_NAND2_NUM843_OUT, XNOR_1_3_NAND2_NUM843_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM843 (.ZN (XNOR_1_1_NAND2_NUM843_OUT), .A1 (N2824), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM843 (.ZN (XNOR_1_2_NAND2_NUM843_OUT), .A1 (GND), .A2 (N1938));
      NOR2_X1 XNOR_1_3_NAND2_NUM843 (.ZN (XNOR_1_3_NAND2_NUM843_OUT), .A1 (XNOR_1_1_NAND2_NUM843_OUT), .A2 (XNOR_1_2_NAND2_NUM843_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM843 (.ZN (N2854), .A1 (XNOR_1_3_NAND2_NUM843_OUT), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM844 (.ZN (N2857), .A1 (N2812), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM845 (.ZN (N2858), .A1 (N2815), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM846 (.ZN (N2859), .A1 (N2818), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM847 (.ZN (N2860), .A1 (N2821), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM848 (.ZN (N2861), .A1 (N2824), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM849 (.ZN (N2862), .A1 (N2829), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM850_OUT, XNOR_1_2_NAND2_NUM850_OUT, XNOR_1_3_NAND2_NUM850_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM850 (.ZN (XNOR_1_1_NAND2_NUM850_OUT), .A1 (N2829), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM850 (.ZN (XNOR_1_2_NAND2_NUM850_OUT), .A1 (GND), .A2 (N1985));
      NOR2_X1 XNOR_1_3_NAND2_NUM850 (.ZN (XNOR_1_3_NAND2_NUM850_OUT), .A1 (XNOR_1_1_NAND2_NUM850_OUT), .A2 (XNOR_1_2_NAND2_NUM850_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM850 (.ZN (N2863), .A1 (XNOR_1_3_NAND2_NUM850_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM851_OUT, XNOR_1_2_NAND2_NUM851_OUT, XNOR_1_3_NAND2_NUM851_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM851 (.ZN (XNOR_1_1_NAND2_NUM851_OUT), .A1 (N2052), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM851 (.ZN (XNOR_1_2_NAND2_NUM851_OUT), .A1 (GND), .A2 (N2857));
      NOR2_X1 XNOR_1_3_NAND2_NUM851 (.ZN (XNOR_1_3_NAND2_NUM851_OUT), .A1 (XNOR_1_1_NAND2_NUM851_OUT), .A2 (XNOR_1_2_NAND2_NUM851_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM851 (.ZN (N2866), .A1 (XNOR_1_3_NAND2_NUM851_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM852_OUT, XNOR_1_2_NAND2_NUM852_OUT, XNOR_1_3_NAND2_NUM852_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM852 (.ZN (XNOR_1_1_NAND2_NUM852_OUT), .A1 (N2055), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM852 (.ZN (XNOR_1_2_NAND2_NUM852_OUT), .A1 (GND), .A2 (N2858));
      NOR2_X1 XNOR_1_3_NAND2_NUM852 (.ZN (XNOR_1_3_NAND2_NUM852_OUT), .A1 (XNOR_1_1_NAND2_NUM852_OUT), .A2 (XNOR_1_2_NAND2_NUM852_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM852 (.ZN (N2867), .A1 (XNOR_1_3_NAND2_NUM852_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM853_OUT, XNOR_1_2_NAND2_NUM853_OUT, XNOR_1_3_NAND2_NUM853_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM853 (.ZN (XNOR_1_1_NAND2_NUM853_OUT), .A1 (N1866), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM853 (.ZN (XNOR_1_2_NAND2_NUM853_OUT), .A1 (GND), .A2 (N2859));
      NOR2_X1 XNOR_1_3_NAND2_NUM853 (.ZN (XNOR_1_3_NAND2_NUM853_OUT), .A1 (XNOR_1_1_NAND2_NUM853_OUT), .A2 (XNOR_1_2_NAND2_NUM853_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM853 (.ZN (N2868), .A1 (XNOR_1_3_NAND2_NUM853_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM854_OUT, XNOR_1_2_NAND2_NUM854_OUT, XNOR_1_3_NAND2_NUM854_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM854 (.ZN (XNOR_1_1_NAND2_NUM854_OUT), .A1 (N1818), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM854 (.ZN (XNOR_1_2_NAND2_NUM854_OUT), .A1 (GND), .A2 (N2860));
      NOR2_X1 XNOR_1_3_NAND2_NUM854 (.ZN (XNOR_1_3_NAND2_NUM854_OUT), .A1 (XNOR_1_1_NAND2_NUM854_OUT), .A2 (XNOR_1_2_NAND2_NUM854_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM854 (.ZN (N2869), .A1 (XNOR_1_3_NAND2_NUM854_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM855_OUT, XNOR_1_2_NAND2_NUM855_OUT, XNOR_1_3_NAND2_NUM855_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM855 (.ZN (XNOR_1_1_NAND2_NUM855_OUT), .A1 (N1902), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM855 (.ZN (XNOR_1_2_NAND2_NUM855_OUT), .A1 (GND), .A2 (N2861));
      NOR2_X1 XNOR_1_3_NAND2_NUM855 (.ZN (XNOR_1_3_NAND2_NUM855_OUT), .A1 (XNOR_1_1_NAND2_NUM855_OUT), .A2 (XNOR_1_2_NAND2_NUM855_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM855 (.ZN (N2870), .A1 (XNOR_1_3_NAND2_NUM855_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM856_OUT, XNOR_1_2_NAND2_NUM856_OUT, XNOR_1_3_NAND2_NUM856_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM856 (.ZN (XNOR_1_1_NAND2_NUM856_OUT), .A1 (N2843), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM856 (.ZN (XNOR_1_2_NAND2_NUM856_OUT), .A1 (GND), .A2 (N886));
      NOR2_X1 XNOR_1_3_NAND2_NUM856 (.ZN (XNOR_1_3_NAND2_NUM856_OUT), .A1 (XNOR_1_1_NAND2_NUM856_OUT), .A2 (XNOR_1_2_NAND2_NUM856_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM856 (.ZN (N2871), .A1 (XNOR_1_3_NAND2_NUM856_OUT), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM857 (.ZN (N2872), .A1 (N2843), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM858_OUT, XNOR_1_2_NAND2_NUM858_OUT, XNOR_1_3_NAND2_NUM858_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM858 (.ZN (XNOR_1_1_NAND2_NUM858_OUT), .A1 (N2846), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM858 (.ZN (XNOR_1_2_NAND2_NUM858_OUT), .A1 (GND), .A2 (N887));
      NOR2_X1 XNOR_1_3_NAND2_NUM858 (.ZN (XNOR_1_3_NAND2_NUM858_OUT), .A1 (XNOR_1_1_NAND2_NUM858_OUT), .A2 (XNOR_1_2_NAND2_NUM858_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM858 (.ZN (N2873), .A1 (XNOR_1_3_NAND2_NUM858_OUT), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM859 (.ZN (N2874), .A1 (N2846), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM860_OUT, XNOR_1_2_NAND2_NUM860_OUT, XNOR_1_3_NAND2_NUM860_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM860 (.ZN (XNOR_1_1_NAND2_NUM860_OUT), .A1 (N1933), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM860 (.ZN (XNOR_1_2_NAND2_NUM860_OUT), .A1 (GND), .A2 (N2862));
      NOR2_X1 XNOR_1_3_NAND2_NUM860 (.ZN (XNOR_1_3_NAND2_NUM860_OUT), .A1 (XNOR_1_1_NAND2_NUM860_OUT), .A2 (XNOR_1_2_NAND2_NUM860_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM860 (.ZN (N2875), .A1 (XNOR_1_3_NAND2_NUM860_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM861_OUT, XNOR_1_2_NAND2_NUM861_OUT, XNOR_1_3_NAND2_NUM861_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM861 (.ZN (XNOR_1_1_NAND2_NUM861_OUT), .A1 (N2866), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM861 (.ZN (XNOR_1_2_NAND2_NUM861_OUT), .A1 (GND), .A2 (N2850));
      NOR2_X1 XNOR_1_3_NAND2_NUM861 (.ZN (XNOR_1_3_NAND2_NUM861_OUT), .A1 (XNOR_1_1_NAND2_NUM861_OUT), .A2 (XNOR_1_2_NAND2_NUM861_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM861 (.ZN (N2876), .A1 (XNOR_1_3_NAND2_NUM861_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM862_OUT, XNOR_1_2_NAND2_NUM862_OUT, XNOR_1_3_NAND2_NUM862_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM862 (.ZN (XNOR_1_1_NAND2_NUM862_OUT), .A1 (N2867), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM862 (.ZN (XNOR_1_2_NAND2_NUM862_OUT), .A1 (GND), .A2 (N2851));
      NOR2_X1 XNOR_1_3_NAND2_NUM862 (.ZN (XNOR_1_3_NAND2_NUM862_OUT), .A1 (XNOR_1_1_NAND2_NUM862_OUT), .A2 (XNOR_1_2_NAND2_NUM862_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM862 (.ZN (N2877), .A1 (XNOR_1_3_NAND2_NUM862_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM863_OUT, XNOR_1_2_NAND2_NUM863_OUT, XNOR_1_3_NAND2_NUM863_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM863 (.ZN (XNOR_1_1_NAND2_NUM863_OUT), .A1 (N2868), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM863 (.ZN (XNOR_1_2_NAND2_NUM863_OUT), .A1 (GND), .A2 (N2852));
      NOR2_X1 XNOR_1_3_NAND2_NUM863 (.ZN (XNOR_1_3_NAND2_NUM863_OUT), .A1 (XNOR_1_1_NAND2_NUM863_OUT), .A2 (XNOR_1_2_NAND2_NUM863_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM863 (.ZN (N2878), .A1 (XNOR_1_3_NAND2_NUM863_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM864_OUT, XNOR_1_2_NAND2_NUM864_OUT, XNOR_1_3_NAND2_NUM864_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM864 (.ZN (XNOR_1_1_NAND2_NUM864_OUT), .A1 (N2869), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM864 (.ZN (XNOR_1_2_NAND2_NUM864_OUT), .A1 (GND), .A2 (N2853));
      NOR2_X1 XNOR_1_3_NAND2_NUM864 (.ZN (XNOR_1_3_NAND2_NUM864_OUT), .A1 (XNOR_1_1_NAND2_NUM864_OUT), .A2 (XNOR_1_2_NAND2_NUM864_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM864 (.ZN (N2879), .A1 (XNOR_1_3_NAND2_NUM864_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM865_OUT, XNOR_1_2_NAND2_NUM865_OUT, XNOR_1_3_NAND2_NUM865_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM865 (.ZN (XNOR_1_1_NAND2_NUM865_OUT), .A1 (N2870), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM865 (.ZN (XNOR_1_2_NAND2_NUM865_OUT), .A1 (GND), .A2 (N2854));
      NOR2_X1 XNOR_1_3_NAND2_NUM865 (.ZN (XNOR_1_3_NAND2_NUM865_OUT), .A1 (XNOR_1_1_NAND2_NUM865_OUT), .A2 (XNOR_1_2_NAND2_NUM865_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM865 (.ZN (N2880), .A1 (XNOR_1_3_NAND2_NUM865_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM866_OUT, XNOR_1_2_NAND2_NUM866_OUT, XNOR_1_3_NAND2_NUM866_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM866 (.ZN (XNOR_1_1_NAND2_NUM866_OUT), .A1 (N682), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM866 (.ZN (XNOR_1_2_NAND2_NUM866_OUT), .A1 (GND), .A2 (N2872));
      NOR2_X1 XNOR_1_3_NAND2_NUM866 (.ZN (XNOR_1_3_NAND2_NUM866_OUT), .A1 (XNOR_1_1_NAND2_NUM866_OUT), .A2 (XNOR_1_2_NAND2_NUM866_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM866 (.ZN (N2881), .A1 (XNOR_1_3_NAND2_NUM866_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM867_OUT, XNOR_1_2_NAND2_NUM867_OUT, XNOR_1_3_NAND2_NUM867_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM867 (.ZN (XNOR_1_1_NAND2_NUM867_OUT), .A1 (N685), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM867 (.ZN (XNOR_1_2_NAND2_NUM867_OUT), .A1 (GND), .A2 (N2874));
      NOR2_X1 XNOR_1_3_NAND2_NUM867 (.ZN (XNOR_1_3_NAND2_NUM867_OUT), .A1 (XNOR_1_1_NAND2_NUM867_OUT), .A2 (XNOR_1_2_NAND2_NUM867_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM867 (.ZN (N2882), .A1 (XNOR_1_3_NAND2_NUM867_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM868_OUT, XNOR_1_2_NAND2_NUM868_OUT, XNOR_1_3_NAND2_NUM868_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM868 (.ZN (XNOR_1_1_NAND2_NUM868_OUT), .A1 (N2875), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM868 (.ZN (XNOR_1_2_NAND2_NUM868_OUT), .A1 (GND), .A2 (N2863));
      NOR2_X1 XNOR_1_3_NAND2_NUM868 (.ZN (XNOR_1_3_NAND2_NUM868_OUT), .A1 (XNOR_1_1_NAND2_NUM868_OUT), .A2 (XNOR_1_2_NAND2_NUM868_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM868 (.ZN (N2883), .A1 (XNOR_1_3_NAND2_NUM868_OUT), .A2 (GND));
      wire XNOR_1_1_AND2_NUM869_OUT, XNOR_1_2_AND2_NUM869_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM869 (.ZN (XNOR_1_1_AND2_NUM869_OUT), .A1 (N2876), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM869 (.ZN (XNOR_1_2_AND2_NUM869_OUT), .A1 (GND), .A2 (N550));
      NOR2_X1 XNOR_1_3_AND2_NUM869 (.ZN (N2886), .A1 (XNOR_1_1_AND2_NUM869_OUT), .A2 (XNOR_1_2_AND2_NUM869_OUT));
      wire XNOR_1_1_AND2_NUM870_OUT, XNOR_1_2_AND2_NUM870_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM870 (.ZN (XNOR_1_1_AND2_NUM870_OUT), .A1 (N551), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM870 (.ZN (XNOR_1_2_AND2_NUM870_OUT), .A1 (GND), .A2 (N2877));
      NOR2_X1 XNOR_1_3_AND2_NUM870 (.ZN (N2887), .A1 (XNOR_1_1_AND2_NUM870_OUT), .A2 (XNOR_1_2_AND2_NUM870_OUT));
      wire XNOR_1_1_AND2_NUM871_OUT, XNOR_1_2_AND2_NUM871_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM871 (.ZN (XNOR_1_1_AND2_NUM871_OUT), .A1 (N553), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM871 (.ZN (XNOR_1_2_AND2_NUM871_OUT), .A1 (GND), .A2 (N2878));
      NOR2_X1 XNOR_1_3_AND2_NUM871 (.ZN (N2888), .A1 (XNOR_1_1_AND2_NUM871_OUT), .A2 (XNOR_1_2_AND2_NUM871_OUT));
      wire XNOR_1_1_AND2_NUM872_OUT, XNOR_1_2_AND2_NUM872_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM872 (.ZN (XNOR_1_1_AND2_NUM872_OUT), .A1 (N2879), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM872 (.ZN (XNOR_1_2_AND2_NUM872_OUT), .A1 (GND), .A2 (N554));
      NOR2_X1 XNOR_1_3_AND2_NUM872 (.ZN (N2889), .A1 (XNOR_1_1_AND2_NUM872_OUT), .A2 (XNOR_1_2_AND2_NUM872_OUT));
      wire XNOR_1_1_AND2_NUM873_OUT, XNOR_1_2_AND2_NUM873_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM873 (.ZN (XNOR_1_1_AND2_NUM873_OUT), .A1 (N555), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM873 (.ZN (XNOR_1_2_AND2_NUM873_OUT), .A1 (GND), .A2 (N2880));
      NOR2_X1 XNOR_1_3_AND2_NUM873 (.ZN (N2890), .A1 (XNOR_1_1_AND2_NUM873_OUT), .A2 (XNOR_1_2_AND2_NUM873_OUT));
      wire XNOR_1_1_NAND2_NUM874_OUT, XNOR_1_2_NAND2_NUM874_OUT, XNOR_1_3_NAND2_NUM874_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM874 (.ZN (XNOR_1_1_NAND2_NUM874_OUT), .A1 (N2871), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM874 (.ZN (XNOR_1_2_NAND2_NUM874_OUT), .A1 (GND), .A2 (N2881));
      NOR2_X1 XNOR_1_3_NAND2_NUM874 (.ZN (XNOR_1_3_NAND2_NUM874_OUT), .A1 (XNOR_1_1_NAND2_NUM874_OUT), .A2 (XNOR_1_2_NAND2_NUM874_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM874 (.ZN (N2891), .A1 (XNOR_1_3_NAND2_NUM874_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM875_OUT, XNOR_1_2_NAND2_NUM875_OUT, XNOR_1_3_NAND2_NUM875_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM875 (.ZN (XNOR_1_1_NAND2_NUM875_OUT), .A1 (N2873), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM875 (.ZN (XNOR_1_2_NAND2_NUM875_OUT), .A1 (GND), .A2 (N2882));
      NOR2_X1 XNOR_1_3_NAND2_NUM875 (.ZN (XNOR_1_3_NAND2_NUM875_OUT), .A1 (XNOR_1_1_NAND2_NUM875_OUT), .A2 (XNOR_1_2_NAND2_NUM875_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM875 (.ZN (N2892), .A1 (XNOR_1_3_NAND2_NUM875_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM876_OUT, XNOR_1_2_NAND2_NUM876_OUT, XNOR_1_3_NAND2_NUM876_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM876 (.ZN (XNOR_1_1_NAND2_NUM876_OUT), .A1 (N2883), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM876 (.ZN (XNOR_1_2_NAND2_NUM876_OUT), .A1 (GND), .A2 (N1461));
      NOR2_X1 XNOR_1_3_NAND2_NUM876 (.ZN (XNOR_1_3_NAND2_NUM876_OUT), .A1 (XNOR_1_1_NAND2_NUM876_OUT), .A2 (XNOR_1_2_NAND2_NUM876_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM876 (.ZN (N2895), .A1 (XNOR_1_3_NAND2_NUM876_OUT), .A2 (GND));
      NOR2_X1 XNOR_NOT1_NUM877 (.ZN (N2896), .A1 (N2883), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM878_OUT, XNOR_1_2_NAND2_NUM878_OUT, XNOR_1_3_NAND2_NUM878_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM878 (.ZN (XNOR_1_1_NAND2_NUM878_OUT), .A1 (N1383), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM878 (.ZN (XNOR_1_2_NAND2_NUM878_OUT), .A1 (GND), .A2 (N2896));
      NOR2_X1 XNOR_1_3_NAND2_NUM878 (.ZN (XNOR_1_3_NAND2_NUM878_OUT), .A1 (XNOR_1_1_NAND2_NUM878_OUT), .A2 (XNOR_1_2_NAND2_NUM878_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM878 (.ZN (N2897), .A1 (XNOR_1_3_NAND2_NUM878_OUT), .A2 (GND));
      wire XNOR_1_1_NAND2_NUM879_OUT, XNOR_1_2_NAND2_NUM879_OUT, XNOR_1_3_NAND2_NUM879_OUT;
      NOR2_X1 XNOR_1_1_NAND2_NUM879 (.ZN (XNOR_1_1_NAND2_NUM879_OUT), .A1 (N2895), .A2 (GND));
      NOR2_X1 XNOR_1_2_NAND2_NUM879 (.ZN (XNOR_1_2_NAND2_NUM879_OUT), .A1 (GND), .A2 (N2897));
      NOR2_X1 XNOR_1_3_NAND2_NUM879 (.ZN (XNOR_1_3_NAND2_NUM879_OUT), .A1 (XNOR_1_1_NAND2_NUM879_OUT), .A2 (XNOR_1_2_NAND2_NUM879_OUT));
      NOR2_X1 XNOR_1_4_NAND2_NUM879 (.ZN (N2898), .A1 (XNOR_1_3_NAND2_NUM879_OUT), .A2 (GND));
      wire XNOR_1_1_AND2_NUM880_OUT, XNOR_1_2_AND2_NUM880_OUT;
      NOR2_X1 XNOR_1_1_AND2_NUM880 (.ZN (XNOR_1_1_AND2_NUM880_OUT), .A1 (N2898), .A2 (GND));
      NOR2_X1 XNOR_1_2_AND2_NUM880 (.ZN (XNOR_1_2_AND2_NUM880_OUT), .A1 (GND), .A2 (N552));
      NOR2_X1 XNOR_1_3_AND2_NUM880 (.ZN (N2899), .A1 (XNOR_1_1_AND2_NUM880_OUT), .A2 (XNOR_1_2_AND2_NUM880_OUT));


      wire XNOR_1_1_N2753_TERMINATION_OUT, XNOR_1_2_N2753_TERMINATION_OUT;
      NOR2_X1 XNOR_1_1_N2753_TERMINATION (.ZN (XNOR_1_1_N2753_TERMINATION_OUT), .A1 (N2753), .A2 (GND));
      NOR2_X1 XNOR_1_2_N2753_TERMINATION (.ZN (N2753_TERMINATION), .A1 (XNOR_1_1_N2753_TERMINATION_OUT), .A2 (XNOR_1_2_N2753_TERMINATION_OUT));

      wire XNOR_1_1_N2754_TERMINATION_OUT, XNOR_1_2_N2754_TERMINATION_OUT;
      NOR2_X1 XNOR_1_1_N2754_TERMINATION (.ZN (XNOR_1_1_N2754_TERMINATION_OUT), .A1 (N2754), .A2 (GND));
      NOR2_X1 XNOR_1_2_N2754_TERMINATION (.ZN (N2754_TERMINATION), .A1 (XNOR_1_1_N2754_TERMINATION_OUT), .A2 (XNOR_1_2_N2754_TERMINATION_OUT));

      wire XNOR_1_1_N2755_TERMINATION_OUT, XNOR_1_2_N2755_TERMINATION_OUT;
      NOR2_X1 XNOR_1_1_N2755_TERMINATION (.ZN (XNOR_1_1_N2755_TERMINATION_OUT), .A1 (N2755), .A2 (GND));
      NOR2_X1 XNOR_1_2_N2755_TERMINATION (.ZN (N2755_TERMINATION), .A1 (XNOR_1_1_N2755_TERMINATION_OUT), .A2 (XNOR_1_2_N2755_TERMINATION_OUT));

      wire XNOR_1_1_N2756_TERMINATION_OUT, XNOR_1_2_N2756_TERMINATION_OUT;
      NOR2_X1 XNOR_1_1_N2756_TERMINATION (.ZN (XNOR_1_1_N2756_TERMINATION_OUT), .A1 (N2756), .A2 (GND));
      NOR2_X1 XNOR_1_2_N2756_TERMINATION (.ZN (N2756_TERMINATION), .A1 (XNOR_1_1_N2756_TERMINATION_OUT), .A2 (XNOR_1_2_N2756_TERMINATION_OUT));

      wire XNOR_1_1_N2762_TERMINATION_OUT, XNOR_1_2_N2762_TERMINATION_OUT;
      NOR2_X1 XNOR_1_1_N2762_TERMINATION (.ZN (XNOR_1_1_N2762_TERMINATION_OUT), .A1 (N2762), .A2 (GND));
      NOR2_X1 XNOR_1_2_N2762_TERMINATION (.ZN (N2762_TERMINATION), .A1 (XNOR_1_1_N2762_TERMINATION_OUT), .A2 (XNOR_1_2_N2762_TERMINATION_OUT));

      wire XNOR_1_1_N2767_TERMINATION_OUT, XNOR_1_2_N2767_TERMINATION_OUT;
      NOR2_X1 XNOR_1_1_N2767_TERMINATION (.ZN (XNOR_1_1_N2767_TERMINATION_OUT), .A1 (N2767), .A2 (GND));
      NOR2_X1 XNOR_1_2_N2767_TERMINATION (.ZN (N2767_TERMINATION), .A1 (XNOR_1_1_N2767_TERMINATION_OUT), .A2 (XNOR_1_2_N2767_TERMINATION_OUT));

      wire XNOR_1_1_N2768_TERMINATION_OUT, XNOR_1_2_N2768_TERMINATION_OUT;
      NOR2_X1 XNOR_1_1_N2768_TERMINATION (.ZN (XNOR_1_1_N2768_TERMINATION_OUT), .A1 (N2768), .A2 (GND));
      NOR2_X1 XNOR_1_2_N2768_TERMINATION (.ZN (N2768_TERMINATION), .A1 (XNOR_1_1_N2768_TERMINATION_OUT), .A2 (XNOR_1_2_N2768_TERMINATION_OUT));

      wire XNOR_1_1_N2779_TERMINATION_OUT, XNOR_1_2_N2779_TERMINATION_OUT;
      NOR2_X1 XNOR_1_1_N2779_TERMINATION (.ZN (XNOR_1_1_N2779_TERMINATION_OUT), .A1 (N2779), .A2 (GND));
      NOR2_X1 XNOR_1_2_N2779_TERMINATION (.ZN (N2779_TERMINATION), .A1 (XNOR_1_1_N2779_TERMINATION_OUT), .A2 (XNOR_1_2_N2779_TERMINATION_OUT));

      wire XNOR_1_1_N2780_TERMINATION_OUT, XNOR_1_2_N2780_TERMINATION_OUT;
      NOR2_X1 XNOR_1_1_N2780_TERMINATION (.ZN (XNOR_1_1_N2780_TERMINATION_OUT), .A1 (N2780), .A2 (GND));
      NOR2_X1 XNOR_1_2_N2780_TERMINATION (.ZN (N2780_TERMINATION), .A1 (XNOR_1_1_N2780_TERMINATION_OUT), .A2 (XNOR_1_2_N2780_TERMINATION_OUT));

      wire XNOR_1_1_N2781_TERMINATION_OUT, XNOR_1_2_N2781_TERMINATION_OUT;
      NOR2_X1 XNOR_1_1_N2781_TERMINATION (.ZN (XNOR_1_1_N2781_TERMINATION_OUT), .A1 (N2781), .A2 (GND));
      NOR2_X1 XNOR_1_2_N2781_TERMINATION (.ZN (N2781_TERMINATION), .A1 (XNOR_1_1_N2781_TERMINATION_OUT), .A2 (XNOR_1_2_N2781_TERMINATION_OUT));

      wire XNOR_1_1_N2782_TERMINATION_OUT, XNOR_1_2_N2782_TERMINATION_OUT;
      NOR2_X1 XNOR_1_1_N2782_TERMINATION (.ZN (XNOR_1_1_N2782_TERMINATION_OUT), .A1 (N2782), .A2 (GND));
      NOR2_X1 XNOR_1_2_N2782_TERMINATION (.ZN (N2782_TERMINATION), .A1 (XNOR_1_1_N2782_TERMINATION_OUT), .A2 (XNOR_1_2_N2782_TERMINATION_OUT));

      wire XNOR_1_1_N2783_TERMINATION_OUT, XNOR_1_2_N2783_TERMINATION_OUT;
      NOR2_X1 XNOR_1_1_N2783_TERMINATION (.ZN (XNOR_1_1_N2783_TERMINATION_OUT), .A1 (N2783), .A2 (GND));
      NOR2_X1 XNOR_1_2_N2783_TERMINATION (.ZN (N2783_TERMINATION), .A1 (XNOR_1_1_N2783_TERMINATION_OUT), .A2 (XNOR_1_2_N2783_TERMINATION_OUT));

      wire XNOR_1_1_N2784_TERMINATION_OUT, XNOR_1_2_N2784_TERMINATION_OUT;
      NOR2_X1 XNOR_1_1_N2784_TERMINATION (.ZN (XNOR_1_1_N2784_TERMINATION_OUT), .A1 (N2784), .A2 (GND));
      NOR2_X1 XNOR_1_2_N2784_TERMINATION (.ZN (N2784_TERMINATION), .A1 (XNOR_1_1_N2784_TERMINATION_OUT), .A2 (XNOR_1_2_N2784_TERMINATION_OUT));

      wire XNOR_1_1_N2785_TERMINATION_OUT, XNOR_1_2_N2785_TERMINATION_OUT;
      NOR2_X1 XNOR_1_1_N2785_TERMINATION (.ZN (XNOR_1_1_N2785_TERMINATION_OUT), .A1 (N2785), .A2 (GND));
      NOR2_X1 XNOR_1_2_N2785_TERMINATION (.ZN (N2785_TERMINATION), .A1 (XNOR_1_1_N2785_TERMINATION_OUT), .A2 (XNOR_1_2_N2785_TERMINATION_OUT));

      wire XNOR_1_1_N2786_TERMINATION_OUT, XNOR_1_2_N2786_TERMINATION_OUT;
      NOR2_X1 XNOR_1_1_N2786_TERMINATION (.ZN (XNOR_1_1_N2786_TERMINATION_OUT), .A1 (N2786), .A2 (GND));
      NOR2_X1 XNOR_1_2_N2786_TERMINATION (.ZN (N2786_TERMINATION), .A1 (XNOR_1_1_N2786_TERMINATION_OUT), .A2 (XNOR_1_2_N2786_TERMINATION_OUT));

      wire XNOR_1_1_N2787_TERMINATION_OUT, XNOR_1_2_N2787_TERMINATION_OUT;
      NOR2_X1 XNOR_1_1_N2787_TERMINATION (.ZN (XNOR_1_1_N2787_TERMINATION_OUT), .A1 (N2787), .A2 (GND));
      NOR2_X1 XNOR_1_2_N2787_TERMINATION (.ZN (N2787_TERMINATION), .A1 (XNOR_1_1_N2787_TERMINATION_OUT), .A2 (XNOR_1_2_N2787_TERMINATION_OUT));

      wire XNOR_1_1_N2811_TERMINATION_OUT, XNOR_1_2_N2811_TERMINATION_OUT;
      NOR2_X1 XNOR_1_1_N2811_TERMINATION (.ZN (XNOR_1_1_N2811_TERMINATION_OUT), .A1 (N2811), .A2 (GND));
      NOR2_X1 XNOR_1_2_N2811_TERMINATION (.ZN (N2811_TERMINATION), .A1 (XNOR_1_1_N2811_TERMINATION_OUT), .A2 (XNOR_1_2_N2811_TERMINATION_OUT));

      wire XNOR_1_1_N2886_TERMINATION_OUT, XNOR_1_2_N2886_TERMINATION_OUT;
      NOR2_X1 XNOR_1_1_N2886_TERMINATION (.ZN (XNOR_1_1_N2886_TERMINATION_OUT), .A1 (N2886), .A2 (GND));
      NOR2_X1 XNOR_1_2_N2886_TERMINATION (.ZN (N2886_TERMINATION), .A1 (XNOR_1_1_N2886_TERMINATION_OUT), .A2 (XNOR_1_2_N2886_TERMINATION_OUT));

      wire XNOR_1_1_N2887_TERMINATION_OUT, XNOR_1_2_N2887_TERMINATION_OUT;
      NOR2_X1 XNOR_1_1_N2887_TERMINATION (.ZN (XNOR_1_1_N2887_TERMINATION_OUT), .A1 (N2887), .A2 (GND));
      NOR2_X1 XNOR_1_2_N2887_TERMINATION (.ZN (N2887_TERMINATION), .A1 (XNOR_1_1_N2887_TERMINATION_OUT), .A2 (XNOR_1_2_N2887_TERMINATION_OUT));

      wire XNOR_1_1_N2888_TERMINATION_OUT, XNOR_1_2_N2888_TERMINATION_OUT;
      NOR2_X1 XNOR_1_1_N2888_TERMINATION (.ZN (XNOR_1_1_N2888_TERMINATION_OUT), .A1 (N2888), .A2 (GND));
      NOR2_X1 XNOR_1_2_N2888_TERMINATION (.ZN (N2888_TERMINATION), .A1 (XNOR_1_1_N2888_TERMINATION_OUT), .A2 (XNOR_1_2_N2888_TERMINATION_OUT));

      wire XNOR_1_1_N2889_TERMINATION_OUT, XNOR_1_2_N2889_TERMINATION_OUT;
      NOR2_X1 XNOR_1_1_N2889_TERMINATION (.ZN (XNOR_1_1_N2889_TERMINATION_OUT), .A1 (N2889), .A2 (GND));
      NOR2_X1 XNOR_1_2_N2889_TERMINATION (.ZN (N2889_TERMINATION), .A1 (XNOR_1_1_N2889_TERMINATION_OUT), .A2 (XNOR_1_2_N2889_TERMINATION_OUT));

      wire XNOR_1_1_N2890_TERMINATION_OUT, XNOR_1_2_N2890_TERMINATION_OUT;
      NOR2_X1 XNOR_1_1_N2890_TERMINATION (.ZN (XNOR_1_1_N2890_TERMINATION_OUT), .A1 (N2890), .A2 (GND));
      NOR2_X1 XNOR_1_2_N2890_TERMINATION (.ZN (N2890_TERMINATION), .A1 (XNOR_1_1_N2890_TERMINATION_OUT), .A2 (XNOR_1_2_N2890_TERMINATION_OUT));

      wire XNOR_1_1_N2891_TERMINATION_OUT, XNOR_1_2_N2891_TERMINATION_OUT;
      NOR2_X1 XNOR_1_1_N2891_TERMINATION (.ZN (XNOR_1_1_N2891_TERMINATION_OUT), .A1 (N2891), .A2 (GND));
      NOR2_X1 XNOR_1_2_N2891_TERMINATION (.ZN (N2891_TERMINATION), .A1 (XNOR_1_1_N2891_TERMINATION_OUT), .A2 (XNOR_1_2_N2891_TERMINATION_OUT));

      wire XNOR_1_1_N2892_TERMINATION_OUT, XNOR_1_2_N2892_TERMINATION_OUT;
      NOR2_X1 XNOR_1_1_N2892_TERMINATION (.ZN (XNOR_1_1_N2892_TERMINATION_OUT), .A1 (N2892), .A2 (GND));
      NOR2_X1 XNOR_1_2_N2892_TERMINATION (.ZN (N2892_TERMINATION), .A1 (XNOR_1_1_N2892_TERMINATION_OUT), .A2 (XNOR_1_2_N2892_TERMINATION_OUT));

      wire XNOR_1_1_N2899_TERMINATION_OUT, XNOR_1_2_N2899_TERMINATION_OUT;
      NOR2_X1 XNOR_1_1_N2899_TERMINATION (.ZN (XNOR_1_1_N2899_TERMINATION_OUT), .A1 (N2899), .A2 (GND));
      NOR2_X1 XNOR_1_2_N2899_TERMINATION (.ZN (N2899_TERMINATION), .A1 (XNOR_1_1_N2899_TERMINATION_OUT), .A2 (XNOR_1_2_N2899_TERMINATION_OUT));


endmodule
module inv_chain (myin, myout);
       input myin;
       output myout;

       wire STAGE0, STAGE1, STAGE2, STAGE3, STAGE4, STAGE5, STAGE6, STAGE7, STAGE8, STAGE9, STAGE10, STAGE11, STAGE12, STAGE13, STAGE14, STAGE15, STAGE16, STAGE17, STAGE18, STAGE19, STAGE20, STAGE21, STAGE22, STAGE23, STAGE24, STAGE25, STAGE26, STAGE27, STAGE28, STAGE29, STAGE30, STAGE31, STAGE32, STAGE33, STAGE34, STAGE35, STAGE36, STAGE37, STAGE38, STAGE39, STAGE40, STAGE41, STAGE42, STAGE43, STAGE44, STAGE45, STAGE46, STAGE47, STAGE48, STAGE49, STAGE50, STAGE51, STAGE52, STAGE53, STAGE54, STAGE55, STAGE56, STAGE57, STAGE58, STAGE59, STAGE60, STAGE61, STAGE62, STAGE63, STAGE64, STAGE65, STAGE66, STAGE67, STAGE68, STAGE69, STAGE70, STAGE71, STAGE72, STAGE73, STAGE74, STAGE75, STAGE76, STAGE77, STAGE78, STAGE79, STAGE80, STAGE81, STAGE82, STAGE83, STAGE84, STAGE85, STAGE86, STAGE87, STAGE88, STAGE89, STAGE90, STAGE91, STAGE92, STAGE93, STAGE94, STAGE95, STAGE96, STAGE97, STAGE98, STAGE99, STAGE100, STAGE101, STAGE102, STAGE103, STAGE104, STAGE105, STAGE106, STAGE107, STAGE108, STAGE109, STAGE110, STAGE111, STAGE112, STAGE113, STAGE114, STAGE115, STAGE116, STAGE117, STAGE118;


       INV_X1 INV0 ( .I (myin), .ZN (STAGE0));
       INV_X1 INV1 ( .I (STAGE0), .ZN (STAGE1));
       INV_X1 INV2 ( .I (STAGE1), .ZN (STAGE2));
       INV_X1 INV3 ( .I (STAGE2), .ZN (STAGE3));
       INV_X1 INV4 ( .I (STAGE3), .ZN (STAGE4));
       INV_X1 INV5 ( .I (STAGE4), .ZN (STAGE5));
       INV_X1 INV6 ( .I (STAGE5), .ZN (STAGE6));
       INV_X1 INV7 ( .I (STAGE6), .ZN (STAGE7));
       INV_X1 INV8 ( .I (STAGE7), .ZN (STAGE8));
       INV_X1 INV9 ( .I (STAGE8), .ZN (STAGE9));
       INV_X1 INV10 ( .I (STAGE9), .ZN (STAGE10));
       INV_X1 INV11 ( .I (STAGE10), .ZN (STAGE11));
       INV_X1 INV12 ( .I (STAGE11), .ZN (STAGE12));
       INV_X1 INV13 ( .I (STAGE12), .ZN (STAGE13));
       INV_X1 INV14 ( .I (STAGE13), .ZN (STAGE14));
       INV_X1 INV15 ( .I (STAGE14), .ZN (STAGE15));
       INV_X1 INV16 ( .I (STAGE15), .ZN (STAGE16));
       INV_X1 INV17 ( .I (STAGE16), .ZN (STAGE17));
       INV_X1 INV18 ( .I (STAGE17), .ZN (STAGE18));
       INV_X1 INV19 ( .I (STAGE18), .ZN (STAGE19));
       INV_X1 INV20 ( .I (STAGE19), .ZN (STAGE20));
       INV_X1 INV21 ( .I (STAGE20), .ZN (STAGE21));
       INV_X1 INV22 ( .I (STAGE21), .ZN (STAGE22));
       INV_X1 INV23 ( .I (STAGE22), .ZN (STAGE23));
       INV_X1 INV24 ( .I (STAGE23), .ZN (STAGE24));
       INV_X1 INV25 ( .I (STAGE24), .ZN (STAGE25));
       INV_X1 INV26 ( .I (STAGE25), .ZN (STAGE26));
       INV_X1 INV27 ( .I (STAGE26), .ZN (STAGE27));
       INV_X1 INV28 ( .I (STAGE27), .ZN (STAGE28));
       INV_X1 INV29 ( .I (STAGE28), .ZN (STAGE29));
       INV_X1 INV30 ( .I (STAGE29), .ZN (STAGE30));
       INV_X1 INV31 ( .I (STAGE30), .ZN (STAGE31));
       INV_X1 INV32 ( .I (STAGE31), .ZN (STAGE32));
       INV_X1 INV33 ( .I (STAGE32), .ZN (STAGE33));
       INV_X1 INV34 ( .I (STAGE33), .ZN (STAGE34));
       INV_X1 INV35 ( .I (STAGE34), .ZN (STAGE35));
       INV_X1 INV36 ( .I (STAGE35), .ZN (STAGE36));
       INV_X1 INV37 ( .I (STAGE36), .ZN (STAGE37));
       INV_X1 INV38 ( .I (STAGE37), .ZN (STAGE38));
       INV_X1 INV39 ( .I (STAGE38), .ZN (STAGE39));
       INV_X1 INV40 ( .I (STAGE39), .ZN (STAGE40));
       INV_X1 INV41 ( .I (STAGE40), .ZN (STAGE41));
       INV_X1 INV42 ( .I (STAGE41), .ZN (STAGE42));
       INV_X1 INV43 ( .I (STAGE42), .ZN (STAGE43));
       INV_X1 INV44 ( .I (STAGE43), .ZN (STAGE44));
       INV_X1 INV45 ( .I (STAGE44), .ZN (STAGE45));
       INV_X1 INV46 ( .I (STAGE45), .ZN (STAGE46));
       INV_X1 INV47 ( .I (STAGE46), .ZN (STAGE47));
       INV_X1 INV48 ( .I (STAGE47), .ZN (STAGE48));
       INV_X1 INV49 ( .I (STAGE48), .ZN (STAGE49));
       INV_X1 INV50 ( .I (STAGE49), .ZN (STAGE50));
       INV_X1 INV51 ( .I (STAGE50), .ZN (STAGE51));
       INV_X1 INV52 ( .I (STAGE51), .ZN (STAGE52));
       INV_X1 INV53 ( .I (STAGE52), .ZN (STAGE53));
       INV_X1 INV54 ( .I (STAGE53), .ZN (STAGE54));
       INV_X1 INV55 ( .I (STAGE54), .ZN (STAGE55));
       INV_X1 INV56 ( .I (STAGE55), .ZN (STAGE56));
       INV_X1 INV57 ( .I (STAGE56), .ZN (STAGE57));
       INV_X1 INV58 ( .I (STAGE57), .ZN (STAGE58));
       INV_X1 INV59 ( .I (STAGE58), .ZN (STAGE59));
       INV_X1 INV60 ( .I (STAGE59), .ZN (STAGE60));
       INV_X1 INV61 ( .I (STAGE60), .ZN (STAGE61));
       INV_X1 INV62 ( .I (STAGE61), .ZN (STAGE62));
       INV_X1 INV63 ( .I (STAGE62), .ZN (STAGE63));
       INV_X1 INV64 ( .I (STAGE63), .ZN (STAGE64));
       INV_X1 INV65 ( .I (STAGE64), .ZN (STAGE65));
       INV_X1 INV66 ( .I (STAGE65), .ZN (STAGE66));
       INV_X1 INV67 ( .I (STAGE66), .ZN (STAGE67));
       INV_X1 INV68 ( .I (STAGE67), .ZN (STAGE68));
       INV_X1 INV69 ( .I (STAGE68), .ZN (STAGE69));
       INV_X1 INV70 ( .I (STAGE69), .ZN (STAGE70));
       INV_X1 INV71 ( .I (STAGE70), .ZN (STAGE71));
       INV_X1 INV72 ( .I (STAGE71), .ZN (STAGE72));
       INV_X1 INV73 ( .I (STAGE72), .ZN (STAGE73));
       INV_X1 INV74 ( .I (STAGE73), .ZN (STAGE74));
       INV_X1 INV75 ( .I (STAGE74), .ZN (STAGE75));
       INV_X1 INV76 ( .I (STAGE75), .ZN (STAGE76));
       INV_X1 INV77 ( .I (STAGE76), .ZN (STAGE77));
       INV_X1 INV78 ( .I (STAGE77), .ZN (STAGE78));
       INV_X1 INV79 ( .I (STAGE78), .ZN (STAGE79));
       INV_X1 INV80 ( .I (STAGE79), .ZN (STAGE80));
       INV_X1 INV81 ( .I (STAGE80), .ZN (STAGE81));
       INV_X1 INV82 ( .I (STAGE81), .ZN (STAGE82));
       INV_X1 INV83 ( .I (STAGE82), .ZN (STAGE83));
       INV_X1 INV84 ( .I (STAGE83), .ZN (STAGE84));
       INV_X1 INV85 ( .I (STAGE84), .ZN (STAGE85));
       INV_X1 INV86 ( .I (STAGE85), .ZN (STAGE86));
       INV_X1 INV87 ( .I (STAGE86), .ZN (STAGE87));
       INV_X1 INV88 ( .I (STAGE87), .ZN (STAGE88));
       INV_X1 INV89 ( .I (STAGE88), .ZN (STAGE89));
       INV_X1 INV90 ( .I (STAGE89), .ZN (STAGE90));
       INV_X1 INV91 ( .I (STAGE90), .ZN (STAGE91));
       INV_X1 INV92 ( .I (STAGE91), .ZN (STAGE92));
       INV_X1 INV93 ( .I (STAGE92), .ZN (STAGE93));
       INV_X1 INV94 ( .I (STAGE93), .ZN (STAGE94));
       INV_X1 INV95 ( .I (STAGE94), .ZN (STAGE95));
       INV_X1 INV96 ( .I (STAGE95), .ZN (STAGE96));
       INV_X1 INV97 ( .I (STAGE96), .ZN (STAGE97));
       INV_X1 INV98 ( .I (STAGE97), .ZN (STAGE98));
       INV_X1 INV99 ( .I (STAGE98), .ZN (STAGE99));
       INV_X1 INV100 ( .I (STAGE99), .ZN (STAGE100));
       INV_X1 INV101 ( .I (STAGE100), .ZN (STAGE101));
       INV_X1 INV102 ( .I (STAGE101), .ZN (STAGE102));
       INV_X1 INV103 ( .I (STAGE102), .ZN (STAGE103));
       INV_X1 INV104 ( .I (STAGE103), .ZN (STAGE104));
       INV_X1 INV105 ( .I (STAGE104), .ZN (STAGE105));
       INV_X1 INV106 ( .I (STAGE105), .ZN (STAGE106));
       INV_X1 INV107 ( .I (STAGE106), .ZN (STAGE107));
       INV_X1 INV108 ( .I (STAGE107), .ZN (STAGE108));
       INV_X1 INV109 ( .I (STAGE108), .ZN (STAGE109));
       INV_X1 INV110 ( .I (STAGE109), .ZN (STAGE110));
       INV_X1 INV111 ( .I (STAGE110), .ZN (STAGE111));
       INV_X1 INV112 ( .I (STAGE111), .ZN (STAGE112));
       INV_X1 INV113 ( .I (STAGE112), .ZN (STAGE113));
       INV_X1 INV114 ( .I (STAGE113), .ZN (STAGE114));
       INV_X1 INV115 ( .I (STAGE114), .ZN (STAGE115));
       INV_X1 INV116 ( .I (STAGE115), .ZN (STAGE116));
       INV_X1 INV117 ( .I (STAGE116), .ZN (STAGE117));
       INV_X1 INV118 ( .I (STAGE117), .ZN (STAGE118));
       INV_X1 INV119 ( .I (STAGE118), .ZN (myout));

endmodule
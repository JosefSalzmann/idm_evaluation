* circuit: nor_A_nor_B_inv_inv_chain
simulator lang=spice

*.PARAM pw=<sed>pw<sed>as
.PARAM supp=0.8V slope=0.1fs
.PARAM t_init0=0.1ns t_init1=0.174ns
.PARAM baseVal=0V peakVal=0.8V tend=1.0ns


.LIB /home/s11777724/involution_tool_library_files/backend/spice/fet.inc CMG

* main circuit
.INCLUDE /home/s11777724/involution_tool_library_files/backend/spice/cell/NOR2_X1.sp
.INCLUDE /home/s11777724/involution_tool_library_files/backend/spice/cell/INV_X1.sp

**** SPECTRE Back Annotation
.option spef='../place_and_route/generic_parasitics.spef'
****

.TEMP 25
.OPTION
+ INGOLD=2
+ PARHIER=LOCAL
*+ POST=CSDF
+ PROBE
+ BRIEF
+ ACCURATE
+ ABSVAR=0.0001
+ DVDT=2
+ RELTOL=1e-11
*+ DELMAX=100fs
+ dc_pivot_check=yes

* vdd
VDD VDD GND 0.8v

VIN myin GND PWL 0ns baseVal t_init0 baseVal 't_init0+slope' peakVal t_init1 peakVal 't_init1+slope' baseVal

* circuit under test
XNOR0 myin GND STAGE0 VDD VDD GND GND NOR2_X1
XNOR1 GND STAGE0 STAGE1 VDD VDD GND GND NOR2_X1
XINV2 STAGE1 STAGE2 VDD VDD GND GND INV_X1

XNOR3 STAGE2 GND STAGE3 VDD VDD GND GND NOR2_X1
XNOR4 GND STAGE3 STAGE4 VDD VDD GND GND NOR2_X1
XINV5 STAGE4 STAGE5 VDD VDD GND GND INV_X1

XNOR6 STAGE5 GND STAGE6 VDD VDD GND GND NOR2_X1
XNOR7 GND STAGE6 STAGE7 VDD VDD GND GND NOR2_X1
XINV8 STAGE7 STAGE8 VDD VDD GND GND INV_X1

XNOR9 STAGE8 GND STAGE9 VDD VDD GND GND NOR2_X1
XNOR10 GND STAGE9 STAGE10 VDD VDD GND GND NOR2_X1
XINV11 STAGE10 STAGE11 VDD VDD GND GND INV_X1

XNOR12 STAGE11 GND STAGE12 VDD VDD GND GND NOR2_X1
XNOR13 GND STAGE12 STAGE13 VDD VDD GND GND NOR2_X1
XINV14 STAGE13 STAGE14 VDD VDD GND GND INV_X1

XNOR15 STAGE14 GND STAGE15 VDD VDD GND GND NOR2_X1
XNOR16 GND STAGE15 STAGE16 VDD VDD GND GND NOR2_X1
XINV17 STAGE16 STAGE17 VDD VDD GND GND INV_X1

XNOR18 STAGE17 GND STAGE18 VDD VDD GND GND NOR2_X1
XNOR19 GND STAGE18 STAGE19 VDD VDD GND GND NOR2_X1
XINV20 STAGE19 STAGE20 VDD VDD GND GND INV_X1

XNOR21 STAGE20 GND STAGE21 VDD VDD GND GND NOR2_X1
XNOR22 GND STAGE21 STAGE22 VDD VDD GND GND NOR2_X1
XINV23 STAGE22 STAGE23 VDD VDD GND GND INV_X1

XNOR24 STAGE23 GND STAGE24 VDD VDD GND GND NOR2_X1
XNOR25 GND STAGE24 STAGE25 VDD VDD GND GND NOR2_X1
XINV26 STAGE25 STAGE26 VDD VDD GND GND INV_X1

XNOR27 STAGE26 GND STAGE27 VDD VDD GND GND NOR2_X1
XNOR28 GND STAGE27 STAGE28 VDD VDD GND GND NOR2_X1
XINV29 STAGE28 STAGE29 VDD VDD GND GND INV_X1

XNOR30 STAGE29 GND STAGE30 VDD VDD GND GND NOR2_X1
XNOR31 GND STAGE30 STAGE31 VDD VDD GND GND NOR2_X1
XINV32 STAGE31 STAGE32 VDD VDD GND GND INV_X1

XNOR33 STAGE32 GND STAGE33 VDD VDD GND GND NOR2_X1
XNOR34 GND STAGE33 STAGE34 VDD VDD GND GND NOR2_X1
XINV35 STAGE34 STAGE35 VDD VDD GND GND INV_X1

XNOR36 STAGE35 GND STAGE36 VDD VDD GND GND NOR2_X1
XNOR37 GND STAGE36 STAGE37 VDD VDD GND GND NOR2_X1
XINV38 STAGE37 O_C_TERM VDD VDD GND GND INV_X1
C_TERM O_C_TERM GND 0.0779pF

.PROBE TRAN V(myin) V(STAGE0) V(STAGE1) V(STAGE2) V(STAGE3) V(STAGE4)
+ V(STAGE5) V(STAGE6) V(STAGE7) V(STAGE8) V(STAGE9) V(STAGE10)
+ V(STAGE11) V(STAGE12) V(STAGE13) V(STAGE14) V(STAGE15)
+ V(STAGE16) V(STAGE17) V(STAGE18) V(STAGE19) V(STAGE20)
+ V(STAGE21) V(STAGE22) V(STAGE23) V(STAGE24) V(STAGE25)
+ V(STAGE26) V(STAGE27) V(STAGE28) V(STAGE29) V(STAGE30)
+ V(STAGE31) V(STAGE32) V(STAGE33) V(STAGE34) V(STAGE35)
+ V(STAGE36) V(STAGE37) V(O_C_TERM)
.TRAN 0.1ps tend
.END
